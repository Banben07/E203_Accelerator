`define TANH_LUT_POSITIVE_SIZE 2140
`define TANH_LUT_POSITIVE_BITS 12
`define TANH_LUT_POSITIVE_0000 16'h0000
`define TANH_LUT_POSITIVE_0008 16'h0008
`define TANH_LUT_POSITIVE_0010 16'h0010
`define TANH_LUT_POSITIVE_0018 16'h0018
`define TANH_LUT_POSITIVE_0020 16'h0020
`define TANH_LUT_POSITIVE_0028 16'h0028
`define TANH_LUT_POSITIVE_0030 16'h0030
`define TANH_LUT_POSITIVE_0038 16'h0038
`define TANH_LUT_POSITIVE_0040 16'h0040
`define TANH_LUT_POSITIVE_0048 16'h0048
`define TANH_LUT_POSITIVE_0050 16'h0050
`define TANH_LUT_POSITIVE_0058 16'h0058
`define TANH_LUT_POSITIVE_0060 16'h0060
`define TANH_LUT_POSITIVE_0068 16'h0068
`define TANH_LUT_POSITIVE_0070 16'h0070
`define TANH_LUT_POSITIVE_0078 16'h0078
`define TANH_LUT_POSITIVE_0080 16'h0080
`define TANH_LUT_POSITIVE_0088 16'h0088
`define TANH_LUT_POSITIVE_0090 16'h0090
`define TANH_LUT_POSITIVE_0098 16'h0098
`define TANH_LUT_POSITIVE_00A0 16'h00A0
`define TANH_LUT_POSITIVE_00A8 16'h00A8
`define TANH_LUT_POSITIVE_00B0 16'h00B0
`define TANH_LUT_POSITIVE_00B8 16'h00B8
`define TANH_LUT_POSITIVE_00C0 16'h00C0
`define TANH_LUT_POSITIVE_00C8 16'h00C8
`define TANH_LUT_POSITIVE_00D0 16'h00D0
`define TANH_LUT_POSITIVE_00D8 16'h00D8
`define TANH_LUT_POSITIVE_00E0 16'h00E0
`define TANH_LUT_POSITIVE_00E8 16'h00E8
`define TANH_LUT_POSITIVE_00F0 16'h00F0
`define TANH_LUT_POSITIVE_00F8 16'h00F8
`define TANH_LUT_POSITIVE_0100 16'h0100
`define TANH_LUT_POSITIVE_0108 16'h0108
`define TANH_LUT_POSITIVE_0110 16'h0110
`define TANH_LUT_POSITIVE_0118 16'h0118
`define TANH_LUT_POSITIVE_0120 16'h0120
`define TANH_LUT_POSITIVE_0128 16'h0128
`define TANH_LUT_POSITIVE_0130 16'h0130
`define TANH_LUT_POSITIVE_0138 16'h0138
`define TANH_LUT_POSITIVE_0140 16'h0140
`define TANH_LUT_POSITIVE_0148 16'h0148
`define TANH_LUT_POSITIVE_0150 16'h0150
`define TANH_LUT_POSITIVE_0158 16'h0158
`define TANH_LUT_POSITIVE_0160 16'h0160
`define TANH_LUT_POSITIVE_0168 16'h0168
`define TANH_LUT_POSITIVE_0170 16'h0170
`define TANH_LUT_POSITIVE_0178 16'h0178
`define TANH_LUT_POSITIVE_0180 16'h0180
`define TANH_LUT_POSITIVE_0188 16'h0188
`define TANH_LUT_POSITIVE_0190 16'h0190
`define TANH_LUT_POSITIVE_0198 16'h0198
`define TANH_LUT_POSITIVE_01A0 16'h01A0
`define TANH_LUT_POSITIVE_01A8 16'h01A8
`define TANH_LUT_POSITIVE_01B0 16'h01B0
`define TANH_LUT_POSITIVE_01B8 16'h01B8
`define TANH_LUT_POSITIVE_01C0 16'h01C0
`define TANH_LUT_POSITIVE_01C8 16'h01C8
`define TANH_LUT_POSITIVE_01D0 16'h01D0
`define TANH_LUT_POSITIVE_01D8 16'h01D8
`define TANH_LUT_POSITIVE_01E0 16'h01E0
`define TANH_LUT_POSITIVE_01E8 16'h01E8
`define TANH_LUT_POSITIVE_01F0 16'h01F0
`define TANH_LUT_POSITIVE_01F8 16'h01F8
`define TANH_LUT_POSITIVE_0200 16'h0200
`define TANH_LUT_POSITIVE_0208 16'h0208
`define TANH_LUT_POSITIVE_0210 16'h0210
`define TANH_LUT_POSITIVE_0218 16'h0218
`define TANH_LUT_POSITIVE_0220 16'h0220
`define TANH_LUT_POSITIVE_0228 16'h0228
`define TANH_LUT_POSITIVE_0230 16'h0230
`define TANH_LUT_POSITIVE_0238 16'h0238
`define TANH_LUT_POSITIVE_0240 16'h0240
`define TANH_LUT_POSITIVE_0248 16'h0248
`define TANH_LUT_POSITIVE_0250 16'h0250
`define TANH_LUT_POSITIVE_0258 16'h0258
`define TANH_LUT_POSITIVE_0260 16'h0260
`define TANH_LUT_POSITIVE_0268 16'h0268
`define TANH_LUT_POSITIVE_0270 16'h0270
`define TANH_LUT_POSITIVE_0278 16'h0278
`define TANH_LUT_POSITIVE_0280 16'h0280
`define TANH_LUT_POSITIVE_0288 16'h0288
`define TANH_LUT_POSITIVE_0290 16'h0290
`define TANH_LUT_POSITIVE_0298 16'h0298
`define TANH_LUT_POSITIVE_02A0 16'h02A0
`define TANH_LUT_POSITIVE_02A8 16'h02A8
`define TANH_LUT_POSITIVE_02B0 16'h02B0
`define TANH_LUT_POSITIVE_02B8 16'h02B8
`define TANH_LUT_POSITIVE_02C0 16'h02C0
`define TANH_LUT_POSITIVE_02C8 16'h02C8
`define TANH_LUT_POSITIVE_02D0 16'h02D0
`define TANH_LUT_POSITIVE_02D8 16'h02D8
`define TANH_LUT_POSITIVE_02E0 16'h02E0
`define TANH_LUT_POSITIVE_02E8 16'h02E8
`define TANH_LUT_POSITIVE_02F0 16'h02F0
`define TANH_LUT_POSITIVE_02F8 16'h02F8
`define TANH_LUT_POSITIVE_0300 16'h0300
`define TANH_LUT_POSITIVE_0308 16'h0308
`define TANH_LUT_POSITIVE_0310 16'h0310
`define TANH_LUT_POSITIVE_0318 16'h0318
`define TANH_LUT_POSITIVE_0320 16'h0320
`define TANH_LUT_POSITIVE_0328 16'h0328
`define TANH_LUT_POSITIVE_0330 16'h0330
`define TANH_LUT_POSITIVE_0338 16'h0338
`define TANH_LUT_POSITIVE_0340 16'h0340
`define TANH_LUT_POSITIVE_0348 16'h0348
`define TANH_LUT_POSITIVE_0350 16'h0350
`define TANH_LUT_POSITIVE_0358 16'h0358
`define TANH_LUT_POSITIVE_0360 16'h0360
`define TANH_LUT_POSITIVE_0368 16'h0368
`define TANH_LUT_POSITIVE_0370 16'h0370
`define TANH_LUT_POSITIVE_0378 16'h0378
`define TANH_LUT_POSITIVE_0380 16'h0380
`define TANH_LUT_POSITIVE_0388 16'h0388
`define TANH_LUT_POSITIVE_0390 16'h0390
`define TANH_LUT_POSITIVE_0398 16'h0398
`define TANH_LUT_POSITIVE_03A0 16'h03A0
`define TANH_LUT_POSITIVE_03A8 16'h03A8
`define TANH_LUT_POSITIVE_03B0 16'h03B0
`define TANH_LUT_POSITIVE_03B8 16'h03B8
`define TANH_LUT_POSITIVE_03C0 16'h03C0
`define TANH_LUT_POSITIVE_03C8 16'h03C8
`define TANH_LUT_POSITIVE_03D0 16'h03D0
`define TANH_LUT_POSITIVE_03D8 16'h03D8
`define TANH_LUT_POSITIVE_03E0 16'h03E0
`define TANH_LUT_POSITIVE_03E8 16'h03E8
`define TANH_LUT_POSITIVE_03F0 16'h03F0
`define TANH_LUT_POSITIVE_03F8 16'h03F8
`define TANH_LUT_POSITIVE_0400 16'h0400
`define TANH_LUT_POSITIVE_0408 16'h0408
`define TANH_LUT_POSITIVE_0410 16'h0410
`define TANH_LUT_POSITIVE_0418 16'h0418
`define TANH_LUT_POSITIVE_0420 16'h0420
`define TANH_LUT_POSITIVE_0428 16'h0428
`define TANH_LUT_POSITIVE_0430 16'h0430
`define TANH_LUT_POSITIVE_0438 16'h0438
`define TANH_LUT_POSITIVE_0440 16'h0440
`define TANH_LUT_POSITIVE_0448 16'h0448
`define TANH_LUT_POSITIVE_0450 16'h0450
`define TANH_LUT_POSITIVE_0458 16'h0458
`define TANH_LUT_POSITIVE_0460 16'h0460
`define TANH_LUT_POSITIVE_0468 16'h0468
`define TANH_LUT_POSITIVE_0470 16'h0470
`define TANH_LUT_POSITIVE_0478 16'h0478
`define TANH_LUT_POSITIVE_0480 16'h0480
`define TANH_LUT_POSITIVE_0488 16'h0488
`define TANH_LUT_POSITIVE_0490 16'h0490
`define TANH_LUT_POSITIVE_0498 16'h0498
`define TANH_LUT_POSITIVE_04A0 16'h04A0
`define TANH_LUT_POSITIVE_04A8 16'h04A8
`define TANH_LUT_POSITIVE_04B0 16'h04B0
`define TANH_LUT_POSITIVE_04B8 16'h04B8
`define TANH_LUT_POSITIVE_04C0 16'h04C0
`define TANH_LUT_POSITIVE_04C8 16'h04C8
`define TANH_LUT_POSITIVE_04D0 16'h04D0
`define TANH_LUT_POSITIVE_04D8 16'h04D8
`define TANH_LUT_POSITIVE_04E0 16'h04E0
`define TANH_LUT_POSITIVE_04E8 16'h04E8
`define TANH_LUT_POSITIVE_04F0 16'h04F0
`define TANH_LUT_POSITIVE_04F8 16'h04F8
`define TANH_LUT_POSITIVE_0500 16'h0500
`define TANH_LUT_POSITIVE_0508 16'h0508
`define TANH_LUT_POSITIVE_0510 16'h0510
`define TANH_LUT_POSITIVE_0518 16'h0518
`define TANH_LUT_POSITIVE_0520 16'h0520
`define TANH_LUT_POSITIVE_0528 16'h0528
`define TANH_LUT_POSITIVE_0530 16'h0530
`define TANH_LUT_POSITIVE_0538 16'h0538
`define TANH_LUT_POSITIVE_0540 16'h0540
`define TANH_LUT_POSITIVE_0548 16'h0548
`define TANH_LUT_POSITIVE_0550 16'h0550
`define TANH_LUT_POSITIVE_0558 16'h0558
`define TANH_LUT_POSITIVE_0560 16'h0560
`define TANH_LUT_POSITIVE_0568 16'h0568
`define TANH_LUT_POSITIVE_0570 16'h0570
`define TANH_LUT_POSITIVE_0578 16'h0578
`define TANH_LUT_POSITIVE_0580 16'h0580
`define TANH_LUT_POSITIVE_0588 16'h0588
`define TANH_LUT_POSITIVE_0590 16'h0590
`define TANH_LUT_POSITIVE_0598 16'h0598
`define TANH_LUT_POSITIVE_05A0 16'h05A0
`define TANH_LUT_POSITIVE_05A8 16'h05A8
`define TANH_LUT_POSITIVE_05B0 16'h05B0
`define TANH_LUT_POSITIVE_05B8 16'h05B8
`define TANH_LUT_POSITIVE_05C0 16'h05C0
`define TANH_LUT_POSITIVE_05C8 16'h05C8
`define TANH_LUT_POSITIVE_05D0 16'h05D0
`define TANH_LUT_POSITIVE_05D8 16'h05D8
`define TANH_LUT_POSITIVE_05E0 16'h05E0
`define TANH_LUT_POSITIVE_05E8 16'h05E8
`define TANH_LUT_POSITIVE_05F0 16'h05F0
`define TANH_LUT_POSITIVE_05F8 16'h05F8
`define TANH_LUT_POSITIVE_0600 16'h0600
`define TANH_LUT_POSITIVE_0608 16'h0608
`define TANH_LUT_POSITIVE_0610 16'h0610
`define TANH_LUT_POSITIVE_0618 16'h0618
`define TANH_LUT_POSITIVE_0620 16'h0620
`define TANH_LUT_POSITIVE_0628 16'h0628
`define TANH_LUT_POSITIVE_0630 16'h0630
`define TANH_LUT_POSITIVE_0638 16'h0638
`define TANH_LUT_POSITIVE_0640 16'h0640
`define TANH_LUT_POSITIVE_0648 16'h0648
`define TANH_LUT_POSITIVE_0650 16'h0650
`define TANH_LUT_POSITIVE_0658 16'h0658
`define TANH_LUT_POSITIVE_0660 16'h0660
`define TANH_LUT_POSITIVE_0668 16'h0668
`define TANH_LUT_POSITIVE_0670 16'h0670
`define TANH_LUT_POSITIVE_0678 16'h0678
`define TANH_LUT_POSITIVE_0680 16'h0680
`define TANH_LUT_POSITIVE_0688 16'h0688
`define TANH_LUT_POSITIVE_0690 16'h0690
`define TANH_LUT_POSITIVE_0698 16'h0698
`define TANH_LUT_POSITIVE_06A0 16'h06A0
`define TANH_LUT_POSITIVE_06A8 16'h06A8
`define TANH_LUT_POSITIVE_06B0 16'h06B0
`define TANH_LUT_POSITIVE_06B8 16'h06B8
`define TANH_LUT_POSITIVE_06C0 16'h06C0
`define TANH_LUT_POSITIVE_06C8 16'h06C8
`define TANH_LUT_POSITIVE_06D0 16'h06D0
`define TANH_LUT_POSITIVE_06D8 16'h06D8
`define TANH_LUT_POSITIVE_06E0 16'h06E0
`define TANH_LUT_POSITIVE_06E8 16'h06E8
`define TANH_LUT_POSITIVE_06F0 16'h06F0
`define TANH_LUT_POSITIVE_06F8 16'h06F8
`define TANH_LUT_POSITIVE_0700 16'h0700
`define TANH_LUT_POSITIVE_0708 16'h0708
`define TANH_LUT_POSITIVE_0710 16'h0710
`define TANH_LUT_POSITIVE_0718 16'h0718
`define TANH_LUT_POSITIVE_0720 16'h0720
`define TANH_LUT_POSITIVE_0728 16'h0728
`define TANH_LUT_POSITIVE_0730 16'h0730
`define TANH_LUT_POSITIVE_0738 16'h0738
`define TANH_LUT_POSITIVE_0740 16'h0740
`define TANH_LUT_POSITIVE_0748 16'h0748
`define TANH_LUT_POSITIVE_0750 16'h0750
`define TANH_LUT_POSITIVE_0758 16'h0758
`define TANH_LUT_POSITIVE_0760 16'h0760
`define TANH_LUT_POSITIVE_0768 16'h0768
`define TANH_LUT_POSITIVE_0770 16'h0770
`define TANH_LUT_POSITIVE_0778 16'h0778
`define TANH_LUT_POSITIVE_0780 16'h0780
`define TANH_LUT_POSITIVE_0788 16'h0788
`define TANH_LUT_POSITIVE_0790 16'h0790
`define TANH_LUT_POSITIVE_0798 16'h0798
`define TANH_LUT_POSITIVE_07A0 16'h07A0
`define TANH_LUT_POSITIVE_07A8 16'h07A8
`define TANH_LUT_POSITIVE_07B0 16'h07B0
`define TANH_LUT_POSITIVE_07B8 16'h07B8
`define TANH_LUT_POSITIVE_07C0 16'h07C0
`define TANH_LUT_POSITIVE_07C8 16'h07C8
`define TANH_LUT_POSITIVE_07D0 16'h07D0
`define TANH_LUT_POSITIVE_07D8 16'h07D8
`define TANH_LUT_POSITIVE_07E0 16'h07E0
`define TANH_LUT_POSITIVE_07E8 16'h07E8
`define TANH_LUT_POSITIVE_07F0 16'h07F0
`define TANH_LUT_POSITIVE_07F8 16'h07F8
`define TANH_LUT_POSITIVE_0800 16'h0800
`define TANH_LUT_POSITIVE_0808 16'h0808
`define TANH_LUT_POSITIVE_0810 16'h0810
`define TANH_LUT_POSITIVE_0818 16'h0818
`define TANH_LUT_POSITIVE_0820 16'h0820
`define TANH_LUT_POSITIVE_0828 16'h0828
`define TANH_LUT_POSITIVE_0830 16'h0830
`define TANH_LUT_POSITIVE_0838 16'h0838
`define TANH_LUT_POSITIVE_0840 16'h0840
`define TANH_LUT_POSITIVE_0848 16'h0848
`define TANH_LUT_POSITIVE_0850 16'h0850
`define TANH_LUT_POSITIVE_0858 16'h0858
`define TANH_LUT_POSITIVE_0860 16'h0860
`define TANH_LUT_POSITIVE_0868 16'h0868
`define TANH_LUT_POSITIVE_0870 16'h0870
`define TANH_LUT_POSITIVE_0878 16'h0878
`define TANH_LUT_POSITIVE_0880 16'h0880
`define TANH_LUT_POSITIVE_0888 16'h0888
`define TANH_LUT_POSITIVE_0890 16'h0890
`define TANH_LUT_POSITIVE_0898 16'h0898
`define TANH_LUT_POSITIVE_08A0 16'h08A0
`define TANH_LUT_POSITIVE_08A8 16'h08A8
`define TANH_LUT_POSITIVE_08B0 16'h08B0
`define TANH_LUT_POSITIVE_08B8 16'h08B8
`define TANH_LUT_POSITIVE_08C0 16'h08C0
`define TANH_LUT_POSITIVE_08C8 16'h08C8
`define TANH_LUT_POSITIVE_08D0 16'h08D0
`define TANH_LUT_POSITIVE_08D8 16'h08D8
`define TANH_LUT_POSITIVE_08E0 16'h08E0
`define TANH_LUT_POSITIVE_08E8 16'h08E8
`define TANH_LUT_POSITIVE_08F0 16'h08F0
`define TANH_LUT_POSITIVE_08F8 16'h08F8
`define TANH_LUT_POSITIVE_0900 16'h0900
`define TANH_LUT_POSITIVE_0908 16'h0908
`define TANH_LUT_POSITIVE_0910 16'h0910
`define TANH_LUT_POSITIVE_0918 16'h0918
`define TANH_LUT_POSITIVE_0920 16'h0920
`define TANH_LUT_POSITIVE_0928 16'h0928
`define TANH_LUT_POSITIVE_0930 16'h0930
`define TANH_LUT_POSITIVE_0938 16'h0938
`define TANH_LUT_POSITIVE_0940 16'h0940
`define TANH_LUT_POSITIVE_0948 16'h0948
`define TANH_LUT_POSITIVE_0950 16'h0950
`define TANH_LUT_POSITIVE_0958 16'h0958
`define TANH_LUT_POSITIVE_0960 16'h0960
`define TANH_LUT_POSITIVE_0968 16'h0968
`define TANH_LUT_POSITIVE_0970 16'h0970
`define TANH_LUT_POSITIVE_0978 16'h0978
`define TANH_LUT_POSITIVE_0980 16'h0980
`define TANH_LUT_POSITIVE_0988 16'h0988
`define TANH_LUT_POSITIVE_0990 16'h0990
`define TANH_LUT_POSITIVE_0998 16'h0998
`define TANH_LUT_POSITIVE_09A0 16'h09A0
`define TANH_LUT_POSITIVE_09A8 16'h09A8
`define TANH_LUT_POSITIVE_09B0 16'h09B0
`define TANH_LUT_POSITIVE_09B8 16'h09B8
`define TANH_LUT_POSITIVE_09C0 16'h09C0
`define TANH_LUT_POSITIVE_09C8 16'h09C8
`define TANH_LUT_POSITIVE_09D0 16'h09D0
`define TANH_LUT_POSITIVE_09D8 16'h09D8
`define TANH_LUT_POSITIVE_09E0 16'h09E0
`define TANH_LUT_POSITIVE_09E8 16'h09E8
`define TANH_LUT_POSITIVE_09F0 16'h09F0
`define TANH_LUT_POSITIVE_09F8 16'h09F8
`define TANH_LUT_POSITIVE_0A00 16'h0A00
`define TANH_LUT_POSITIVE_0A08 16'h0A08
`define TANH_LUT_POSITIVE_0A10 16'h0A10
`define TANH_LUT_POSITIVE_0A18 16'h0A18
`define TANH_LUT_POSITIVE_0A20 16'h0A20
`define TANH_LUT_POSITIVE_0A28 16'h0A28
`define TANH_LUT_POSITIVE_0A30 16'h0A30
`define TANH_LUT_POSITIVE_0A38 16'h0A38
`define TANH_LUT_POSITIVE_0A40 16'h0A40
`define TANH_LUT_POSITIVE_0A48 16'h0A48
`define TANH_LUT_POSITIVE_0A50 16'h0A50
`define TANH_LUT_POSITIVE_0A58 16'h0A58
`define TANH_LUT_POSITIVE_0A60 16'h0A60
`define TANH_LUT_POSITIVE_0A68 16'h0A68
`define TANH_LUT_POSITIVE_0A70 16'h0A70
`define TANH_LUT_POSITIVE_0A78 16'h0A78
`define TANH_LUT_POSITIVE_0A80 16'h0A80
`define TANH_LUT_POSITIVE_0A88 16'h0A88
`define TANH_LUT_POSITIVE_0A90 16'h0A90
`define TANH_LUT_POSITIVE_0A98 16'h0A98
`define TANH_LUT_POSITIVE_0AA0 16'h0AA0
`define TANH_LUT_POSITIVE_0AA8 16'h0AA8
`define TANH_LUT_POSITIVE_0AB0 16'h0AB0
`define TANH_LUT_POSITIVE_0AB8 16'h0AB8
`define TANH_LUT_POSITIVE_0AC0 16'h0AC0
`define TANH_LUT_POSITIVE_0AC8 16'h0AC8
`define TANH_LUT_POSITIVE_0AD0 16'h0AD0
`define TANH_LUT_POSITIVE_0AD8 16'h0AD8
`define TANH_LUT_POSITIVE_0AE0 16'h0AE0
`define TANH_LUT_POSITIVE_0AE8 16'h0AE8
`define TANH_LUT_POSITIVE_0AF0 16'h0AF0
`define TANH_LUT_POSITIVE_0AF8 16'h0AF8
`define TANH_LUT_POSITIVE_0B00 16'h0B00
`define TANH_LUT_POSITIVE_0B08 16'h0B08
`define TANH_LUT_POSITIVE_0B10 16'h0B10
`define TANH_LUT_POSITIVE_0B18 16'h0B18
`define TANH_LUT_POSITIVE_0B20 16'h0B20
`define TANH_LUT_POSITIVE_0B28 16'h0B28
`define TANH_LUT_POSITIVE_0B30 16'h0B30
`define TANH_LUT_POSITIVE_0B38 16'h0B38
`define TANH_LUT_POSITIVE_0B40 16'h0B40
`define TANH_LUT_POSITIVE_0B48 16'h0B48
`define TANH_LUT_POSITIVE_0B50 16'h0B50
`define TANH_LUT_POSITIVE_0B58 16'h0B58
`define TANH_LUT_POSITIVE_0B60 16'h0B60
`define TANH_LUT_POSITIVE_0B68 16'h0B68
`define TANH_LUT_POSITIVE_0B70 16'h0B70
`define TANH_LUT_POSITIVE_0B78 16'h0B78
`define TANH_LUT_POSITIVE_0B80 16'h0B80
`define TANH_LUT_POSITIVE_0B88 16'h0B88
`define TANH_LUT_POSITIVE_0B90 16'h0B90
`define TANH_LUT_POSITIVE_0B98 16'h0B98
`define TANH_LUT_POSITIVE_0BA0 16'h0BA0
`define TANH_LUT_POSITIVE_0BA8 16'h0BA8
`define TANH_LUT_POSITIVE_0BB0 16'h0BB0
`define TANH_LUT_POSITIVE_0BB8 16'h0BB8
`define TANH_LUT_POSITIVE_0BC0 16'h0BC0
`define TANH_LUT_POSITIVE_0BC8 16'h0BC8
`define TANH_LUT_POSITIVE_0BD0 16'h0BD0
`define TANH_LUT_POSITIVE_0BD8 16'h0BD8
`define TANH_LUT_POSITIVE_0BE0 16'h0BE0
`define TANH_LUT_POSITIVE_0BE8 16'h0BE8
`define TANH_LUT_POSITIVE_0BF0 16'h0BF0
`define TANH_LUT_POSITIVE_0BF8 16'h0BF8
`define TANH_LUT_POSITIVE_0C00 16'h0C00
`define TANH_LUT_POSITIVE_0C08 16'h0C08
`define TANH_LUT_POSITIVE_0C10 16'h0C10
`define TANH_LUT_POSITIVE_0C18 16'h0C18
`define TANH_LUT_POSITIVE_0C20 16'h0C20
`define TANH_LUT_POSITIVE_0C28 16'h0C28
`define TANH_LUT_POSITIVE_0C30 16'h0C30
`define TANH_LUT_POSITIVE_0C38 16'h0C38
`define TANH_LUT_POSITIVE_0C40 16'h0C40
`define TANH_LUT_POSITIVE_0C48 16'h0C48
`define TANH_LUT_POSITIVE_0C50 16'h0C50
`define TANH_LUT_POSITIVE_0C58 16'h0C58
`define TANH_LUT_POSITIVE_0C60 16'h0C60
`define TANH_LUT_POSITIVE_0C68 16'h0C68
`define TANH_LUT_POSITIVE_0C70 16'h0C70
`define TANH_LUT_POSITIVE_0C78 16'h0C78
`define TANH_LUT_POSITIVE_0C80 16'h0C80
`define TANH_LUT_POSITIVE_0C88 16'h0C88
`define TANH_LUT_POSITIVE_0C90 16'h0C90
`define TANH_LUT_POSITIVE_0C98 16'h0C98
`define TANH_LUT_POSITIVE_0CA0 16'h0CA0
`define TANH_LUT_POSITIVE_0CA8 16'h0CA8
`define TANH_LUT_POSITIVE_0CB0 16'h0CB0
`define TANH_LUT_POSITIVE_0CB8 16'h0CB8
`define TANH_LUT_POSITIVE_0CC0 16'h0CC0
`define TANH_LUT_POSITIVE_0CC8 16'h0CC8
`define TANH_LUT_POSITIVE_0CD0 16'h0CD0
`define TANH_LUT_POSITIVE_0CD8 16'h0CD8
`define TANH_LUT_POSITIVE_0CE0 16'h0CE0
`define TANH_LUT_POSITIVE_0CE8 16'h0CE8
`define TANH_LUT_POSITIVE_0CF0 16'h0CF0
`define TANH_LUT_POSITIVE_0CF8 16'h0CF8
`define TANH_LUT_POSITIVE_0D00 16'h0D00
`define TANH_LUT_POSITIVE_0D08 16'h0D08
`define TANH_LUT_POSITIVE_0D10 16'h0D10
`define TANH_LUT_POSITIVE_0D18 16'h0D18
`define TANH_LUT_POSITIVE_0D20 16'h0D20
`define TANH_LUT_POSITIVE_0D28 16'h0D28
`define TANH_LUT_POSITIVE_0D30 16'h0D30
`define TANH_LUT_POSITIVE_0D38 16'h0D38
`define TANH_LUT_POSITIVE_0D40 16'h0D40
`define TANH_LUT_POSITIVE_0D48 16'h0D48
`define TANH_LUT_POSITIVE_0D50 16'h0D50
`define TANH_LUT_POSITIVE_0D58 16'h0D58
`define TANH_LUT_POSITIVE_0D60 16'h0D60
`define TANH_LUT_POSITIVE_0D68 16'h0D68
`define TANH_LUT_POSITIVE_0D70 16'h0D70
`define TANH_LUT_POSITIVE_0D78 16'h0D78
`define TANH_LUT_POSITIVE_0D80 16'h0D80
`define TANH_LUT_POSITIVE_0D88 16'h0D88
`define TANH_LUT_POSITIVE_0D90 16'h0D90
`define TANH_LUT_POSITIVE_0D98 16'h0D98
`define TANH_LUT_POSITIVE_0DA0 16'h0DA0
`define TANH_LUT_POSITIVE_0DA8 16'h0DA8
`define TANH_LUT_POSITIVE_0DB0 16'h0DB0
`define TANH_LUT_POSITIVE_0DB8 16'h0DB8
`define TANH_LUT_POSITIVE_0DC0 16'h0DC0
`define TANH_LUT_POSITIVE_0DC8 16'h0DC8
`define TANH_LUT_POSITIVE_0DD0 16'h0DD0
`define TANH_LUT_POSITIVE_0DD8 16'h0DD8
`define TANH_LUT_POSITIVE_0DE0 16'h0DE0
`define TANH_LUT_POSITIVE_0DE8 16'h0DE8
`define TANH_LUT_POSITIVE_0DF0 16'h0DF0
`define TANH_LUT_POSITIVE_0DF8 16'h0DF8
`define TANH_LUT_POSITIVE_0E00 16'h0E00
`define TANH_LUT_POSITIVE_0E08 16'h0E08
`define TANH_LUT_POSITIVE_0E10 16'h0E10
`define TANH_LUT_POSITIVE_0E18 16'h0E18
`define TANH_LUT_POSITIVE_0E20 16'h0E20
`define TANH_LUT_POSITIVE_0E28 16'h0E28
`define TANH_LUT_POSITIVE_0E30 16'h0E30
`define TANH_LUT_POSITIVE_0E38 16'h0E38
`define TANH_LUT_POSITIVE_0E40 16'h0E40
`define TANH_LUT_POSITIVE_0E48 16'h0E48
`define TANH_LUT_POSITIVE_0E50 16'h0E50
`define TANH_LUT_POSITIVE_0E58 16'h0E58
`define TANH_LUT_POSITIVE_0E60 16'h0E60
`define TANH_LUT_POSITIVE_0E68 16'h0E68
`define TANH_LUT_POSITIVE_0E70 16'h0E70
`define TANH_LUT_POSITIVE_0E78 16'h0E78
`define TANH_LUT_POSITIVE_0E80 16'h0E80
`define TANH_LUT_POSITIVE_0E88 16'h0E88
`define TANH_LUT_POSITIVE_0E90 16'h0E90
`define TANH_LUT_POSITIVE_0E98 16'h0E98
`define TANH_LUT_POSITIVE_0EA0 16'h0EA0
`define TANH_LUT_POSITIVE_0EA8 16'h0EA8
`define TANH_LUT_POSITIVE_0EB0 16'h0EB0
`define TANH_LUT_POSITIVE_0EB8 16'h0EB8
`define TANH_LUT_POSITIVE_0EC0 16'h0EC0
`define TANH_LUT_POSITIVE_0EC8 16'h0EC8
`define TANH_LUT_POSITIVE_0ED0 16'h0ED0
`define TANH_LUT_POSITIVE_0ED8 16'h0ED8
`define TANH_LUT_POSITIVE_0EE0 16'h0EE0
`define TANH_LUT_POSITIVE_0EE8 16'h0EE8
`define TANH_LUT_POSITIVE_0EF0 16'h0EF0
`define TANH_LUT_POSITIVE_0EF8 16'h0EF8
`define TANH_LUT_POSITIVE_0F00 16'h0F00
`define TANH_LUT_POSITIVE_0F08 16'h0F08
`define TANH_LUT_POSITIVE_0F10 16'h0F10
`define TANH_LUT_POSITIVE_0F18 16'h0F18
`define TANH_LUT_POSITIVE_0F20 16'h0F20
`define TANH_LUT_POSITIVE_0F28 16'h0F28
`define TANH_LUT_POSITIVE_0F30 16'h0F30
`define TANH_LUT_POSITIVE_0F38 16'h0F38
`define TANH_LUT_POSITIVE_0F40 16'h0F40
`define TANH_LUT_POSITIVE_0F48 16'h0F48
`define TANH_LUT_POSITIVE_0F50 16'h0F50
`define TANH_LUT_POSITIVE_0F58 16'h0F58
`define TANH_LUT_POSITIVE_0F60 16'h0F60
`define TANH_LUT_POSITIVE_0F68 16'h0F68
`define TANH_LUT_POSITIVE_0F70 16'h0F70
`define TANH_LUT_POSITIVE_0F78 16'h0F78
`define TANH_LUT_POSITIVE_0F80 16'h0F80
`define TANH_LUT_POSITIVE_0F88 16'h0F88
`define TANH_LUT_POSITIVE_0F90 16'h0F90
`define TANH_LUT_POSITIVE_0F98 16'h0F98
`define TANH_LUT_POSITIVE_0FA0 16'h0FA0
`define TANH_LUT_POSITIVE_0FA8 16'h0FA8
`define TANH_LUT_POSITIVE_0FB0 16'h0FB0
`define TANH_LUT_POSITIVE_0FB8 16'h0FB8
`define TANH_LUT_POSITIVE_0FC0 16'h0FC0
`define TANH_LUT_POSITIVE_0FC8 16'h0FC8
`define TANH_LUT_POSITIVE_0FD0 16'h0FD0
`define TANH_LUT_POSITIVE_0FD8 16'h0FD8
`define TANH_LUT_POSITIVE_0FE0 16'h0FE0
`define TANH_LUT_POSITIVE_0FE8 16'h0FE8
`define TANH_LUT_POSITIVE_0FF0 16'h0FF0
`define TANH_LUT_POSITIVE_0FF8 16'h0FF8
`define TANH_LUT_POSITIVE_1000 16'h1000
`define TANH_LUT_POSITIVE_1008 16'h1008
`define TANH_LUT_POSITIVE_1010 16'h1010
`define TANH_LUT_POSITIVE_1018 16'h1018
`define TANH_LUT_POSITIVE_1020 16'h1020
`define TANH_LUT_POSITIVE_1028 16'h1028
`define TANH_LUT_POSITIVE_1030 16'h1030
`define TANH_LUT_POSITIVE_1038 16'h1038
`define TANH_LUT_POSITIVE_1040 16'h1040
`define TANH_LUT_POSITIVE_1048 16'h1048
`define TANH_LUT_POSITIVE_1050 16'h1050
`define TANH_LUT_POSITIVE_1058 16'h1058
`define TANH_LUT_POSITIVE_1060 16'h1060
`define TANH_LUT_POSITIVE_1068 16'h1068
`define TANH_LUT_POSITIVE_1070 16'h1070
`define TANH_LUT_POSITIVE_1078 16'h1078
`define TANH_LUT_POSITIVE_1080 16'h1080
`define TANH_LUT_POSITIVE_1088 16'h1088
`define TANH_LUT_POSITIVE_1090 16'h1090
`define TANH_LUT_POSITIVE_1098 16'h1098
`define TANH_LUT_POSITIVE_10A0 16'h10A0
`define TANH_LUT_POSITIVE_10A8 16'h10A8
`define TANH_LUT_POSITIVE_10B0 16'h10B0
`define TANH_LUT_POSITIVE_10B8 16'h10B8
`define TANH_LUT_POSITIVE_10C0 16'h10C0
`define TANH_LUT_POSITIVE_10C8 16'h10C8
`define TANH_LUT_POSITIVE_10D0 16'h10D0
`define TANH_LUT_POSITIVE_10D8 16'h10D8
`define TANH_LUT_POSITIVE_10E0 16'h10E0
`define TANH_LUT_POSITIVE_10E8 16'h10E8
`define TANH_LUT_POSITIVE_10F0 16'h10F0
`define TANH_LUT_POSITIVE_10F8 16'h10F8
`define TANH_LUT_POSITIVE_1100 16'h1100
`define TANH_LUT_POSITIVE_1108 16'h1108
`define TANH_LUT_POSITIVE_1110 16'h1110
`define TANH_LUT_POSITIVE_1118 16'h1118
`define TANH_LUT_POSITIVE_1120 16'h1120
`define TANH_LUT_POSITIVE_1128 16'h1128
`define TANH_LUT_POSITIVE_1130 16'h1130
`define TANH_LUT_POSITIVE_1138 16'h1138
`define TANH_LUT_POSITIVE_1140 16'h1140
`define TANH_LUT_POSITIVE_1148 16'h1148
`define TANH_LUT_POSITIVE_1150 16'h1150
`define TANH_LUT_POSITIVE_1158 16'h1158
`define TANH_LUT_POSITIVE_1160 16'h1160
`define TANH_LUT_POSITIVE_1168 16'h1168
`define TANH_LUT_POSITIVE_1170 16'h1170
`define TANH_LUT_POSITIVE_1178 16'h1178
`define TANH_LUT_POSITIVE_1180 16'h1180
`define TANH_LUT_POSITIVE_1188 16'h1188
`define TANH_LUT_POSITIVE_1190 16'h1190
`define TANH_LUT_POSITIVE_1198 16'h1198
`define TANH_LUT_POSITIVE_11A0 16'h11A0
`define TANH_LUT_POSITIVE_11A8 16'h11A8
`define TANH_LUT_POSITIVE_11B0 16'h11B0
`define TANH_LUT_POSITIVE_11B8 16'h11B8
`define TANH_LUT_POSITIVE_11C0 16'h11C0
`define TANH_LUT_POSITIVE_11C8 16'h11C8
`define TANH_LUT_POSITIVE_11D0 16'h11D0
`define TANH_LUT_POSITIVE_11D8 16'h11D8
`define TANH_LUT_POSITIVE_11E0 16'h11E0
`define TANH_LUT_POSITIVE_11E8 16'h11E8
`define TANH_LUT_POSITIVE_11F0 16'h11F0
`define TANH_LUT_POSITIVE_11F8 16'h11F8
`define TANH_LUT_POSITIVE_1200 16'h1200
`define TANH_LUT_POSITIVE_1208 16'h1208
`define TANH_LUT_POSITIVE_1210 16'h1210
`define TANH_LUT_POSITIVE_1218 16'h1218
`define TANH_LUT_POSITIVE_1220 16'h1220
`define TANH_LUT_POSITIVE_1228 16'h1228
`define TANH_LUT_POSITIVE_1230 16'h1230
`define TANH_LUT_POSITIVE_1238 16'h1238
`define TANH_LUT_POSITIVE_1240 16'h1240
`define TANH_LUT_POSITIVE_1248 16'h1248
`define TANH_LUT_POSITIVE_1250 16'h1250
`define TANH_LUT_POSITIVE_1258 16'h1258
`define TANH_LUT_POSITIVE_1260 16'h1260
`define TANH_LUT_POSITIVE_1268 16'h1268
`define TANH_LUT_POSITIVE_1270 16'h1270
`define TANH_LUT_POSITIVE_1278 16'h1278
`define TANH_LUT_POSITIVE_1280 16'h1280
`define TANH_LUT_POSITIVE_1288 16'h1288
`define TANH_LUT_POSITIVE_1290 16'h1290
`define TANH_LUT_POSITIVE_1298 16'h1298
`define TANH_LUT_POSITIVE_12A0 16'h12A0
`define TANH_LUT_POSITIVE_12A8 16'h12A8
`define TANH_LUT_POSITIVE_12B0 16'h12B0
`define TANH_LUT_POSITIVE_12B8 16'h12B8
`define TANH_LUT_POSITIVE_12C0 16'h12C0
`define TANH_LUT_POSITIVE_12C8 16'h12C8
`define TANH_LUT_POSITIVE_12D0 16'h12D0
`define TANH_LUT_POSITIVE_12D8 16'h12D8
`define TANH_LUT_POSITIVE_12E0 16'h12E0
`define TANH_LUT_POSITIVE_12E8 16'h12E8
`define TANH_LUT_POSITIVE_12F0 16'h12F0
`define TANH_LUT_POSITIVE_12F8 16'h12F8
`define TANH_LUT_POSITIVE_1300 16'h1300
`define TANH_LUT_POSITIVE_1308 16'h1308
`define TANH_LUT_POSITIVE_1310 16'h1310
`define TANH_LUT_POSITIVE_1318 16'h1318
`define TANH_LUT_POSITIVE_1320 16'h1320
`define TANH_LUT_POSITIVE_1328 16'h1328
`define TANH_LUT_POSITIVE_1330 16'h1330
`define TANH_LUT_POSITIVE_1338 16'h1338
`define TANH_LUT_POSITIVE_1340 16'h1340
`define TANH_LUT_POSITIVE_1348 16'h1348
`define TANH_LUT_POSITIVE_1350 16'h1350
`define TANH_LUT_POSITIVE_1358 16'h1358
`define TANH_LUT_POSITIVE_1360 16'h1360
`define TANH_LUT_POSITIVE_1368 16'h1368
`define TANH_LUT_POSITIVE_1370 16'h1370
`define TANH_LUT_POSITIVE_1378 16'h1378
`define TANH_LUT_POSITIVE_1380 16'h1380
`define TANH_LUT_POSITIVE_1388 16'h1388
`define TANH_LUT_POSITIVE_1390 16'h1390
`define TANH_LUT_POSITIVE_1398 16'h1398
`define TANH_LUT_POSITIVE_13A0 16'h13A0
`define TANH_LUT_POSITIVE_13A8 16'h13A8
`define TANH_LUT_POSITIVE_13B0 16'h13B0
`define TANH_LUT_POSITIVE_13B8 16'h13B8
`define TANH_LUT_POSITIVE_13C0 16'h13C0
`define TANH_LUT_POSITIVE_13C8 16'h13C8
`define TANH_LUT_POSITIVE_13D0 16'h13D0
`define TANH_LUT_POSITIVE_13D8 16'h13D8
`define TANH_LUT_POSITIVE_13E0 16'h13E0
`define TANH_LUT_POSITIVE_13E8 16'h13E8
`define TANH_LUT_POSITIVE_13F0 16'h13F0
`define TANH_LUT_POSITIVE_13F8 16'h13F8
`define TANH_LUT_POSITIVE_1400 16'h1400
`define TANH_LUT_POSITIVE_1408 16'h1408
`define TANH_LUT_POSITIVE_1410 16'h1410
`define TANH_LUT_POSITIVE_1418 16'h1418
`define TANH_LUT_POSITIVE_1420 16'h1420
`define TANH_LUT_POSITIVE_1428 16'h1428
`define TANH_LUT_POSITIVE_1430 16'h1430
`define TANH_LUT_POSITIVE_1438 16'h1438
`define TANH_LUT_POSITIVE_1440 16'h1440
`define TANH_LUT_POSITIVE_1448 16'h1448
`define TANH_LUT_POSITIVE_1450 16'h1450
`define TANH_LUT_POSITIVE_1458 16'h1458
`define TANH_LUT_POSITIVE_1460 16'h1460
`define TANH_LUT_POSITIVE_1468 16'h1468
`define TANH_LUT_POSITIVE_1470 16'h1470
`define TANH_LUT_POSITIVE_1478 16'h1478
`define TANH_LUT_POSITIVE_1480 16'h1480
`define TANH_LUT_POSITIVE_1488 16'h1488
`define TANH_LUT_POSITIVE_1490 16'h1490
`define TANH_LUT_POSITIVE_1498 16'h1498
`define TANH_LUT_POSITIVE_14A0 16'h14A0
`define TANH_LUT_POSITIVE_14A8 16'h14A8
`define TANH_LUT_POSITIVE_14B0 16'h14B0
`define TANH_LUT_POSITIVE_14B8 16'h14B8
`define TANH_LUT_POSITIVE_14C0 16'h14C0
`define TANH_LUT_POSITIVE_14C8 16'h14C8
`define TANH_LUT_POSITIVE_14D0 16'h14D0
`define TANH_LUT_POSITIVE_14D8 16'h14D8
`define TANH_LUT_POSITIVE_14E0 16'h14E0
`define TANH_LUT_POSITIVE_14E8 16'h14E8
`define TANH_LUT_POSITIVE_14F0 16'h14F0
`define TANH_LUT_POSITIVE_14F8 16'h14F8
`define TANH_LUT_POSITIVE_1500 16'h1500
`define TANH_LUT_POSITIVE_1508 16'h1508
`define TANH_LUT_POSITIVE_1510 16'h1510
`define TANH_LUT_POSITIVE_1518 16'h1518
`define TANH_LUT_POSITIVE_1520 16'h1520
`define TANH_LUT_POSITIVE_1528 16'h1528
`define TANH_LUT_POSITIVE_1530 16'h1530
`define TANH_LUT_POSITIVE_1538 16'h1538
`define TANH_LUT_POSITIVE_1540 16'h1540
`define TANH_LUT_POSITIVE_1548 16'h1548
`define TANH_LUT_POSITIVE_1550 16'h1550
`define TANH_LUT_POSITIVE_1558 16'h1558
`define TANH_LUT_POSITIVE_1560 16'h1560
`define TANH_LUT_POSITIVE_1568 16'h1568
`define TANH_LUT_POSITIVE_1570 16'h1570
`define TANH_LUT_POSITIVE_1578 16'h1578
`define TANH_LUT_POSITIVE_1580 16'h1580
`define TANH_LUT_POSITIVE_1588 16'h1588
`define TANH_LUT_POSITIVE_1590 16'h1590
`define TANH_LUT_POSITIVE_1598 16'h1598
`define TANH_LUT_POSITIVE_15A0 16'h15A0
`define TANH_LUT_POSITIVE_15A8 16'h15A8
`define TANH_LUT_POSITIVE_15B0 16'h15B0
`define TANH_LUT_POSITIVE_15B8 16'h15B8
`define TANH_LUT_POSITIVE_15C0 16'h15C0
`define TANH_LUT_POSITIVE_15C8 16'h15C8
`define TANH_LUT_POSITIVE_15D0 16'h15D0
`define TANH_LUT_POSITIVE_15D8 16'h15D8
`define TANH_LUT_POSITIVE_15E0 16'h15E0
`define TANH_LUT_POSITIVE_15E8 16'h15E8
`define TANH_LUT_POSITIVE_15F0 16'h15F0
`define TANH_LUT_POSITIVE_15F8 16'h15F8
`define TANH_LUT_POSITIVE_1600 16'h1600
`define TANH_LUT_POSITIVE_1608 16'h1608
`define TANH_LUT_POSITIVE_1610 16'h1610
`define TANH_LUT_POSITIVE_1618 16'h1618
`define TANH_LUT_POSITIVE_1620 16'h1620
`define TANH_LUT_POSITIVE_1628 16'h1628
`define TANH_LUT_POSITIVE_1630 16'h1630
`define TANH_LUT_POSITIVE_1638 16'h1638
`define TANH_LUT_POSITIVE_1640 16'h1640
`define TANH_LUT_POSITIVE_1648 16'h1648
`define TANH_LUT_POSITIVE_1650 16'h1650
`define TANH_LUT_POSITIVE_1658 16'h1658
`define TANH_LUT_POSITIVE_1660 16'h1660
`define TANH_LUT_POSITIVE_1668 16'h1668
`define TANH_LUT_POSITIVE_1670 16'h1670
`define TANH_LUT_POSITIVE_1678 16'h1678
`define TANH_LUT_POSITIVE_1680 16'h1680
`define TANH_LUT_POSITIVE_1688 16'h1688
`define TANH_LUT_POSITIVE_1690 16'h1690
`define TANH_LUT_POSITIVE_1698 16'h1698
`define TANH_LUT_POSITIVE_16A0 16'h16A0
`define TANH_LUT_POSITIVE_16A8 16'h16A8
`define TANH_LUT_POSITIVE_16B0 16'h16B0
`define TANH_LUT_POSITIVE_16B8 16'h16B8
`define TANH_LUT_POSITIVE_16C0 16'h16C0
`define TANH_LUT_POSITIVE_16C8 16'h16C8
`define TANH_LUT_POSITIVE_16D0 16'h16D0
`define TANH_LUT_POSITIVE_16D8 16'h16D8
`define TANH_LUT_POSITIVE_16E0 16'h16E0
`define TANH_LUT_POSITIVE_16E8 16'h16E8
`define TANH_LUT_POSITIVE_16F0 16'h16F0
`define TANH_LUT_POSITIVE_16F8 16'h16F8
`define TANH_LUT_POSITIVE_1700 16'h1700
`define TANH_LUT_POSITIVE_1708 16'h1708
`define TANH_LUT_POSITIVE_1710 16'h1710
`define TANH_LUT_POSITIVE_1718 16'h1718
`define TANH_LUT_POSITIVE_1720 16'h1720
`define TANH_LUT_POSITIVE_1728 16'h1728
`define TANH_LUT_POSITIVE_1730 16'h1730
`define TANH_LUT_POSITIVE_1738 16'h1738
`define TANH_LUT_POSITIVE_1740 16'h1740
`define TANH_LUT_POSITIVE_1748 16'h1748
`define TANH_LUT_POSITIVE_1750 16'h1750
`define TANH_LUT_POSITIVE_1758 16'h1758
`define TANH_LUT_POSITIVE_1760 16'h1760
`define TANH_LUT_POSITIVE_1768 16'h1768
`define TANH_LUT_POSITIVE_1770 16'h1770
`define TANH_LUT_POSITIVE_1778 16'h1778
`define TANH_LUT_POSITIVE_1780 16'h1780
`define TANH_LUT_POSITIVE_1788 16'h1788
`define TANH_LUT_POSITIVE_1790 16'h1790
`define TANH_LUT_POSITIVE_1798 16'h1798
`define TANH_LUT_POSITIVE_17A0 16'h17A0
`define TANH_LUT_POSITIVE_17A8 16'h17A8
`define TANH_LUT_POSITIVE_17B0 16'h17B0
`define TANH_LUT_POSITIVE_17B8 16'h17B8
`define TANH_LUT_POSITIVE_17C0 16'h17C0
`define TANH_LUT_POSITIVE_17C8 16'h17C8
`define TANH_LUT_POSITIVE_17D0 16'h17D0
`define TANH_LUT_POSITIVE_17D8 16'h17D8
`define TANH_LUT_POSITIVE_17E0 16'h17E0
`define TANH_LUT_POSITIVE_17E8 16'h17E8
`define TANH_LUT_POSITIVE_17F0 16'h17F0
`define TANH_LUT_POSITIVE_17F8 16'h17F8
`define TANH_LUT_POSITIVE_1800 16'h1800
`define TANH_LUT_POSITIVE_1808 16'h1808
`define TANH_LUT_POSITIVE_1810 16'h1810
`define TANH_LUT_POSITIVE_1818 16'h1818
`define TANH_LUT_POSITIVE_1820 16'h1820
`define TANH_LUT_POSITIVE_1828 16'h1828
`define TANH_LUT_POSITIVE_1830 16'h1830
`define TANH_LUT_POSITIVE_1838 16'h1838
`define TANH_LUT_POSITIVE_1840 16'h1840
`define TANH_LUT_POSITIVE_1848 16'h1848
`define TANH_LUT_POSITIVE_1850 16'h1850
`define TANH_LUT_POSITIVE_1858 16'h1858
`define TANH_LUT_POSITIVE_1860 16'h1860
`define TANH_LUT_POSITIVE_1868 16'h1868
`define TANH_LUT_POSITIVE_1870 16'h1870
`define TANH_LUT_POSITIVE_1878 16'h1878
`define TANH_LUT_POSITIVE_1880 16'h1880
`define TANH_LUT_POSITIVE_1888 16'h1888
`define TANH_LUT_POSITIVE_1890 16'h1890
`define TANH_LUT_POSITIVE_1898 16'h1898
`define TANH_LUT_POSITIVE_18A0 16'h18A0
`define TANH_LUT_POSITIVE_18A8 16'h18A8
`define TANH_LUT_POSITIVE_18B0 16'h18B0
`define TANH_LUT_POSITIVE_18B8 16'h18B8
`define TANH_LUT_POSITIVE_18C0 16'h18C0
`define TANH_LUT_POSITIVE_18C8 16'h18C8
`define TANH_LUT_POSITIVE_18D0 16'h18D0
`define TANH_LUT_POSITIVE_18D8 16'h18D8
`define TANH_LUT_POSITIVE_18E0 16'h18E0
`define TANH_LUT_POSITIVE_18E8 16'h18E8
`define TANH_LUT_POSITIVE_18F0 16'h18F0
`define TANH_LUT_POSITIVE_18F8 16'h18F8
`define TANH_LUT_POSITIVE_1900 16'h1900
`define TANH_LUT_POSITIVE_1908 16'h1908
`define TANH_LUT_POSITIVE_1910 16'h1910
`define TANH_LUT_POSITIVE_1918 16'h1918
`define TANH_LUT_POSITIVE_1920 16'h1920
`define TANH_LUT_POSITIVE_1928 16'h1928
`define TANH_LUT_POSITIVE_1930 16'h1930
`define TANH_LUT_POSITIVE_1938 16'h1938
`define TANH_LUT_POSITIVE_1940 16'h1940
`define TANH_LUT_POSITIVE_1948 16'h1948
`define TANH_LUT_POSITIVE_1950 16'h1950
`define TANH_LUT_POSITIVE_1958 16'h1958
`define TANH_LUT_POSITIVE_1960 16'h1960
`define TANH_LUT_POSITIVE_1968 16'h1968
`define TANH_LUT_POSITIVE_1970 16'h1970
`define TANH_LUT_POSITIVE_1978 16'h1978
`define TANH_LUT_POSITIVE_1980 16'h1980
`define TANH_LUT_POSITIVE_1988 16'h1988
`define TANH_LUT_POSITIVE_1990 16'h1990
`define TANH_LUT_POSITIVE_1998 16'h1998
`define TANH_LUT_POSITIVE_19A0 16'h19A0
`define TANH_LUT_POSITIVE_19A8 16'h19A8
`define TANH_LUT_POSITIVE_19B0 16'h19B0
`define TANH_LUT_POSITIVE_19B8 16'h19B8
`define TANH_LUT_POSITIVE_19C0 16'h19C0
`define TANH_LUT_POSITIVE_19C8 16'h19C8
`define TANH_LUT_POSITIVE_19D0 16'h19D0
`define TANH_LUT_POSITIVE_19D8 16'h19D8
`define TANH_LUT_POSITIVE_19E0 16'h19E0
`define TANH_LUT_POSITIVE_19E8 16'h19E8
`define TANH_LUT_POSITIVE_19F0 16'h19F0
`define TANH_LUT_POSITIVE_19F8 16'h19F8
`define TANH_LUT_POSITIVE_1A00 16'h1A00
`define TANH_LUT_POSITIVE_1A08 16'h1A08
`define TANH_LUT_POSITIVE_1A10 16'h1A10
`define TANH_LUT_POSITIVE_1A18 16'h1A18
`define TANH_LUT_POSITIVE_1A20 16'h1A20
`define TANH_LUT_POSITIVE_1A28 16'h1A28
`define TANH_LUT_POSITIVE_1A30 16'h1A30
`define TANH_LUT_POSITIVE_1A38 16'h1A38
`define TANH_LUT_POSITIVE_1A40 16'h1A40
`define TANH_LUT_POSITIVE_1A48 16'h1A48
`define TANH_LUT_POSITIVE_1A50 16'h1A50
`define TANH_LUT_POSITIVE_1A58 16'h1A58
`define TANH_LUT_POSITIVE_1A60 16'h1A60
`define TANH_LUT_POSITIVE_1A68 16'h1A68
`define TANH_LUT_POSITIVE_1A70 16'h1A70
`define TANH_LUT_POSITIVE_1A78 16'h1A78
`define TANH_LUT_POSITIVE_1A80 16'h1A80
`define TANH_LUT_POSITIVE_1A88 16'h1A88
`define TANH_LUT_POSITIVE_1A90 16'h1A90
`define TANH_LUT_POSITIVE_1A98 16'h1A98
`define TANH_LUT_POSITIVE_1AA0 16'h1AA0
`define TANH_LUT_POSITIVE_1AA8 16'h1AA8
`define TANH_LUT_POSITIVE_1AB0 16'h1AB0
`define TANH_LUT_POSITIVE_1AB8 16'h1AB8
`define TANH_LUT_POSITIVE_1AC0 16'h1AC0
`define TANH_LUT_POSITIVE_1AC8 16'h1AC8
`define TANH_LUT_POSITIVE_1AD0 16'h1AD0
`define TANH_LUT_POSITIVE_1AD8 16'h1AD8
`define TANH_LUT_POSITIVE_1AE0 16'h1AE0
`define TANH_LUT_POSITIVE_1AE8 16'h1AE8
`define TANH_LUT_POSITIVE_1AF0 16'h1AF0
`define TANH_LUT_POSITIVE_1AF8 16'h1AF8
`define TANH_LUT_POSITIVE_1B00 16'h1B00
`define TANH_LUT_POSITIVE_1B08 16'h1B08
`define TANH_LUT_POSITIVE_1B10 16'h1B10
`define TANH_LUT_POSITIVE_1B18 16'h1B18
`define TANH_LUT_POSITIVE_1B20 16'h1B20
`define TANH_LUT_POSITIVE_1B28 16'h1B28
`define TANH_LUT_POSITIVE_1B30 16'h1B30
`define TANH_LUT_POSITIVE_1B38 16'h1B38
`define TANH_LUT_POSITIVE_1B40 16'h1B40
`define TANH_LUT_POSITIVE_1B48 16'h1B48
`define TANH_LUT_POSITIVE_1B50 16'h1B50
`define TANH_LUT_POSITIVE_1B58 16'h1B58
`define TANH_LUT_POSITIVE_1B60 16'h1B60
`define TANH_LUT_POSITIVE_1B68 16'h1B68
`define TANH_LUT_POSITIVE_1B70 16'h1B70
`define TANH_LUT_POSITIVE_1B78 16'h1B78
`define TANH_LUT_POSITIVE_1B80 16'h1B80
`define TANH_LUT_POSITIVE_1B88 16'h1B88
`define TANH_LUT_POSITIVE_1B90 16'h1B90
`define TANH_LUT_POSITIVE_1B98 16'h1B98
`define TANH_LUT_POSITIVE_1BA0 16'h1BA0
`define TANH_LUT_POSITIVE_1BA8 16'h1BA8
`define TANH_LUT_POSITIVE_1BB0 16'h1BB0
`define TANH_LUT_POSITIVE_1BB8 16'h1BB8
`define TANH_LUT_POSITIVE_1BC0 16'h1BC0
`define TANH_LUT_POSITIVE_1BC8 16'h1BC8
`define TANH_LUT_POSITIVE_1BD0 16'h1BD0
`define TANH_LUT_POSITIVE_1BD8 16'h1BD8
`define TANH_LUT_POSITIVE_1BE0 16'h1BE0
`define TANH_LUT_POSITIVE_1BE8 16'h1BE8
`define TANH_LUT_POSITIVE_1BF0 16'h1BF0
`define TANH_LUT_POSITIVE_1BF8 16'h1BF8
`define TANH_LUT_POSITIVE_1C00 16'h1C00
`define TANH_LUT_POSITIVE_1C08 16'h1C08
`define TANH_LUT_POSITIVE_1C10 16'h1C10
`define TANH_LUT_POSITIVE_1C18 16'h1C18
`define TANH_LUT_POSITIVE_1C20 16'h1C20
`define TANH_LUT_POSITIVE_1C28 16'h1C28
`define TANH_LUT_POSITIVE_1C30 16'h1C30
`define TANH_LUT_POSITIVE_1C38 16'h1C38
`define TANH_LUT_POSITIVE_1C40 16'h1C40
`define TANH_LUT_POSITIVE_1C48 16'h1C48
`define TANH_LUT_POSITIVE_1C50 16'h1C50
`define TANH_LUT_POSITIVE_1C58 16'h1C58
`define TANH_LUT_POSITIVE_1C60 16'h1C60
`define TANH_LUT_POSITIVE_1C68 16'h1C68
`define TANH_LUT_POSITIVE_1C70 16'h1C70
`define TANH_LUT_POSITIVE_1C78 16'h1C78
`define TANH_LUT_POSITIVE_1C80 16'h1C80
`define TANH_LUT_POSITIVE_1C88 16'h1C88
`define TANH_LUT_POSITIVE_1C90 16'h1C90
`define TANH_LUT_POSITIVE_1C98 16'h1C98
`define TANH_LUT_POSITIVE_1CA0 16'h1CA0
`define TANH_LUT_POSITIVE_1CA8 16'h1CA8
`define TANH_LUT_POSITIVE_1CB0 16'h1CB0
`define TANH_LUT_POSITIVE_1CB8 16'h1CB8
`define TANH_LUT_POSITIVE_1CC0 16'h1CC0
`define TANH_LUT_POSITIVE_1CC8 16'h1CC8
`define TANH_LUT_POSITIVE_1CD0 16'h1CD0
`define TANH_LUT_POSITIVE_1CD8 16'h1CD8
`define TANH_LUT_POSITIVE_1CE0 16'h1CE0
`define TANH_LUT_POSITIVE_1CE8 16'h1CE8
`define TANH_LUT_POSITIVE_1CF0 16'h1CF0
`define TANH_LUT_POSITIVE_1CF8 16'h1CF8
`define TANH_LUT_POSITIVE_1D00 16'h1D00
`define TANH_LUT_POSITIVE_1D08 16'h1D08
`define TANH_LUT_POSITIVE_1D10 16'h1D10
`define TANH_LUT_POSITIVE_1D18 16'h1D18
`define TANH_LUT_POSITIVE_1D20 16'h1D20
`define TANH_LUT_POSITIVE_1D28 16'h1D28
`define TANH_LUT_POSITIVE_1D30 16'h1D30
`define TANH_LUT_POSITIVE_1D38 16'h1D38
`define TANH_LUT_POSITIVE_1D40 16'h1D40
`define TANH_LUT_POSITIVE_1D48 16'h1D48
`define TANH_LUT_POSITIVE_1D50 16'h1D50
`define TANH_LUT_POSITIVE_1D58 16'h1D58
`define TANH_LUT_POSITIVE_1D60 16'h1D60
`define TANH_LUT_POSITIVE_1D68 16'h1D68
`define TANH_LUT_POSITIVE_1D70 16'h1D70
`define TANH_LUT_POSITIVE_1D78 16'h1D78
`define TANH_LUT_POSITIVE_1D80 16'h1D80
`define TANH_LUT_POSITIVE_1D88 16'h1D88
`define TANH_LUT_POSITIVE_1D90 16'h1D90
`define TANH_LUT_POSITIVE_1D98 16'h1D98
`define TANH_LUT_POSITIVE_1DA0 16'h1DA0
`define TANH_LUT_POSITIVE_1DA8 16'h1DA8
`define TANH_LUT_POSITIVE_1DB0 16'h1DB0
`define TANH_LUT_POSITIVE_1DB8 16'h1DB8
`define TANH_LUT_POSITIVE_1DC0 16'h1DC0
`define TANH_LUT_POSITIVE_1DC8 16'h1DC8
`define TANH_LUT_POSITIVE_1DD0 16'h1DD0
`define TANH_LUT_POSITIVE_1DD8 16'h1DD8
`define TANH_LUT_POSITIVE_1DE0 16'h1DE0
`define TANH_LUT_POSITIVE_1DE8 16'h1DE8
`define TANH_LUT_POSITIVE_1DF0 16'h1DF0
`define TANH_LUT_POSITIVE_1DF8 16'h1DF8
`define TANH_LUT_POSITIVE_1E00 16'h1E00
`define TANH_LUT_POSITIVE_1E08 16'h1E08
`define TANH_LUT_POSITIVE_1E10 16'h1E10
`define TANH_LUT_POSITIVE_1E18 16'h1E18
`define TANH_LUT_POSITIVE_1E20 16'h1E20
`define TANH_LUT_POSITIVE_1E28 16'h1E28
`define TANH_LUT_POSITIVE_1E30 16'h1E30
`define TANH_LUT_POSITIVE_1E38 16'h1E38
`define TANH_LUT_POSITIVE_1E40 16'h1E40
`define TANH_LUT_POSITIVE_1E48 16'h1E48
`define TANH_LUT_POSITIVE_1E50 16'h1E50
`define TANH_LUT_POSITIVE_1E58 16'h1E58
`define TANH_LUT_POSITIVE_1E60 16'h1E60
`define TANH_LUT_POSITIVE_1E68 16'h1E68
`define TANH_LUT_POSITIVE_1E70 16'h1E70
`define TANH_LUT_POSITIVE_1E78 16'h1E78
`define TANH_LUT_POSITIVE_1E80 16'h1E80
`define TANH_LUT_POSITIVE_1E88 16'h1E88
`define TANH_LUT_POSITIVE_1E90 16'h1E90
`define TANH_LUT_POSITIVE_1E98 16'h1E98
`define TANH_LUT_POSITIVE_1EA0 16'h1EA0
`define TANH_LUT_POSITIVE_1EA8 16'h1EA8
`define TANH_LUT_POSITIVE_1EB0 16'h1EB0
`define TANH_LUT_POSITIVE_1EB8 16'h1EB8
`define TANH_LUT_POSITIVE_1EC0 16'h1EC0
`define TANH_LUT_POSITIVE_1EC8 16'h1EC8
`define TANH_LUT_POSITIVE_1ED0 16'h1ED0
`define TANH_LUT_POSITIVE_1ED8 16'h1ED8
`define TANH_LUT_POSITIVE_1EE0 16'h1EE0
`define TANH_LUT_POSITIVE_1EE8 16'h1EE8
`define TANH_LUT_POSITIVE_1EF0 16'h1EF0
`define TANH_LUT_POSITIVE_1EF8 16'h1EF8
`define TANH_LUT_POSITIVE_1F00 16'h1F00
`define TANH_LUT_POSITIVE_1F08 16'h1F08
`define TANH_LUT_POSITIVE_1F10 16'h1F10
`define TANH_LUT_POSITIVE_1F18 16'h1F18
`define TANH_LUT_POSITIVE_1F20 16'h1F20
`define TANH_LUT_POSITIVE_1F28 16'h1F28
`define TANH_LUT_POSITIVE_1F30 16'h1F30
`define TANH_LUT_POSITIVE_1F38 16'h1F38
`define TANH_LUT_POSITIVE_1F40 16'h1F40
`define TANH_LUT_POSITIVE_1F48 16'h1F48
`define TANH_LUT_POSITIVE_1F50 16'h1F50
`define TANH_LUT_POSITIVE_1F58 16'h1F58
`define TANH_LUT_POSITIVE_1F60 16'h1F60
`define TANH_LUT_POSITIVE_1F68 16'h1F68
`define TANH_LUT_POSITIVE_1F70 16'h1F70
`define TANH_LUT_POSITIVE_1F78 16'h1F78
`define TANH_LUT_POSITIVE_1F80 16'h1F80
`define TANH_LUT_POSITIVE_1F88 16'h1F88
`define TANH_LUT_POSITIVE_1F90 16'h1F90
`define TANH_LUT_POSITIVE_1F98 16'h1F98
`define TANH_LUT_POSITIVE_1FA0 16'h1FA0
`define TANH_LUT_POSITIVE_1FA8 16'h1FA8
`define TANH_LUT_POSITIVE_1FB0 16'h1FB0
`define TANH_LUT_POSITIVE_1FB8 16'h1FB8
`define TANH_LUT_POSITIVE_1FC0 16'h1FC0
`define TANH_LUT_POSITIVE_1FC8 16'h1FC8
`define TANH_LUT_POSITIVE_1FD0 16'h1FD0
`define TANH_LUT_POSITIVE_1FD8 16'h1FD8
`define TANH_LUT_POSITIVE_1FE0 16'h1FE0
`define TANH_LUT_POSITIVE_1FE8 16'h1FE8
`define TANH_LUT_POSITIVE_1FF0 16'h1FF0
`define TANH_LUT_POSITIVE_1FF8 16'h1FF8
`define TANH_LUT_POSITIVE_2000 16'h2000
`define TANH_LUT_POSITIVE_2008 16'h2008
`define TANH_LUT_POSITIVE_2010 16'h2010
`define TANH_LUT_POSITIVE_2018 16'h2018
`define TANH_LUT_POSITIVE_2020 16'h2020
`define TANH_LUT_POSITIVE_2028 16'h2028
`define TANH_LUT_POSITIVE_2030 16'h2030
`define TANH_LUT_POSITIVE_2038 16'h2038
`define TANH_LUT_POSITIVE_2040 16'h2040
`define TANH_LUT_POSITIVE_2048 16'h2048
`define TANH_LUT_POSITIVE_2050 16'h2050
`define TANH_LUT_POSITIVE_2058 16'h2058
`define TANH_LUT_POSITIVE_2060 16'h2060
`define TANH_LUT_POSITIVE_2068 16'h2068
`define TANH_LUT_POSITIVE_2070 16'h2070
`define TANH_LUT_POSITIVE_2078 16'h2078
`define TANH_LUT_POSITIVE_2080 16'h2080
`define TANH_LUT_POSITIVE_2088 16'h2088
`define TANH_LUT_POSITIVE_2090 16'h2090
`define TANH_LUT_POSITIVE_2098 16'h2098
`define TANH_LUT_POSITIVE_20A0 16'h20A0
`define TANH_LUT_POSITIVE_20A8 16'h20A8
`define TANH_LUT_POSITIVE_20B0 16'h20B0
`define TANH_LUT_POSITIVE_20B8 16'h20B8
`define TANH_LUT_POSITIVE_20C0 16'h20C0
`define TANH_LUT_POSITIVE_20C8 16'h20C8
`define TANH_LUT_POSITIVE_20D0 16'h20D0
`define TANH_LUT_POSITIVE_20D8 16'h20D8
`define TANH_LUT_POSITIVE_20E0 16'h20E0
`define TANH_LUT_POSITIVE_20E8 16'h20E8
`define TANH_LUT_POSITIVE_20F0 16'h20F0
`define TANH_LUT_POSITIVE_20F8 16'h20F8
`define TANH_LUT_POSITIVE_2100 16'h2100
`define TANH_LUT_POSITIVE_2108 16'h2108
`define TANH_LUT_POSITIVE_2110 16'h2110
`define TANH_LUT_POSITIVE_2118 16'h2118
`define TANH_LUT_POSITIVE_2120 16'h2120
`define TANH_LUT_POSITIVE_2128 16'h2128
`define TANH_LUT_POSITIVE_2130 16'h2130
`define TANH_LUT_POSITIVE_2138 16'h2138
`define TANH_LUT_POSITIVE_2140 16'h2140
`define TANH_LUT_POSITIVE_2148 16'h2148
`define TANH_LUT_POSITIVE_2150 16'h2150
`define TANH_LUT_POSITIVE_2158 16'h2158
`define TANH_LUT_POSITIVE_2160 16'h2160
`define TANH_LUT_POSITIVE_2168 16'h2168
`define TANH_LUT_POSITIVE_2170 16'h2170
`define TANH_LUT_POSITIVE_2178 16'h2178
`define TANH_LUT_POSITIVE_2180 16'h2180
`define TANH_LUT_POSITIVE_2188 16'h2188
`define TANH_LUT_POSITIVE_2190 16'h2190
`define TANH_LUT_POSITIVE_2198 16'h2198
`define TANH_LUT_POSITIVE_21A0 16'h21A0
`define TANH_LUT_POSITIVE_21A8 16'h21A8
`define TANH_LUT_POSITIVE_21B0 16'h21B0
`define TANH_LUT_POSITIVE_21B8 16'h21B8
`define TANH_LUT_POSITIVE_21C0 16'h21C0
`define TANH_LUT_POSITIVE_21C8 16'h21C8
`define TANH_LUT_POSITIVE_21D0 16'h21D0
`define TANH_LUT_POSITIVE_21D8 16'h21D8
`define TANH_LUT_POSITIVE_21E0 16'h21E0
`define TANH_LUT_POSITIVE_21E8 16'h21E8
`define TANH_LUT_POSITIVE_21F0 16'h21F0
`define TANH_LUT_POSITIVE_21F8 16'h21F8
`define TANH_LUT_POSITIVE_2200 16'h2200
`define TANH_LUT_POSITIVE_2208 16'h2208
`define TANH_LUT_POSITIVE_2210 16'h2210
`define TANH_LUT_POSITIVE_2218 16'h2218
`define TANH_LUT_POSITIVE_2220 16'h2220
`define TANH_LUT_POSITIVE_2228 16'h2228
`define TANH_LUT_POSITIVE_2230 16'h2230
`define TANH_LUT_POSITIVE_2238 16'h2238
`define TANH_LUT_POSITIVE_2240 16'h2240
`define TANH_LUT_POSITIVE_2248 16'h2248
`define TANH_LUT_POSITIVE_2250 16'h2250
`define TANH_LUT_POSITIVE_2258 16'h2258
`define TANH_LUT_POSITIVE_2260 16'h2260
`define TANH_LUT_POSITIVE_2268 16'h2268
`define TANH_LUT_POSITIVE_2270 16'h2270
`define TANH_LUT_POSITIVE_2278 16'h2278
`define TANH_LUT_POSITIVE_2280 16'h2280
`define TANH_LUT_POSITIVE_2288 16'h2288
`define TANH_LUT_POSITIVE_2290 16'h2290
`define TANH_LUT_POSITIVE_2298 16'h2298
`define TANH_LUT_POSITIVE_22A0 16'h22A0
`define TANH_LUT_POSITIVE_22A8 16'h22A8
`define TANH_LUT_POSITIVE_22B0 16'h22B0
`define TANH_LUT_POSITIVE_22B8 16'h22B8
`define TANH_LUT_POSITIVE_22C0 16'h22C0
`define TANH_LUT_POSITIVE_22C8 16'h22C8
`define TANH_LUT_POSITIVE_22D0 16'h22D0
`define TANH_LUT_POSITIVE_22D8 16'h22D8
`define TANH_LUT_POSITIVE_22E0 16'h22E0
`define TANH_LUT_POSITIVE_22E8 16'h22E8
`define TANH_LUT_POSITIVE_22F0 16'h22F0
`define TANH_LUT_POSITIVE_22F8 16'h22F8
`define TANH_LUT_POSITIVE_2300 16'h2300
`define TANH_LUT_POSITIVE_2308 16'h2308
`define TANH_LUT_POSITIVE_2310 16'h2310
`define TANH_LUT_POSITIVE_2318 16'h2318
`define TANH_LUT_POSITIVE_2320 16'h2320
`define TANH_LUT_POSITIVE_2328 16'h2328
`define TANH_LUT_POSITIVE_2330 16'h2330
`define TANH_LUT_POSITIVE_2338 16'h2338
`define TANH_LUT_POSITIVE_2340 16'h2340
`define TANH_LUT_POSITIVE_2348 16'h2348
`define TANH_LUT_POSITIVE_2350 16'h2350
`define TANH_LUT_POSITIVE_2358 16'h2358
`define TANH_LUT_POSITIVE_2360 16'h2360
`define TANH_LUT_POSITIVE_2368 16'h2368
`define TANH_LUT_POSITIVE_2370 16'h2370
`define TANH_LUT_POSITIVE_2378 16'h2378
`define TANH_LUT_POSITIVE_2380 16'h2380
`define TANH_LUT_POSITIVE_2388 16'h2388
`define TANH_LUT_POSITIVE_2390 16'h2390
`define TANH_LUT_POSITIVE_2398 16'h2398
`define TANH_LUT_POSITIVE_23A0 16'h23A0
`define TANH_LUT_POSITIVE_23A8 16'h23A8
`define TANH_LUT_POSITIVE_23B0 16'h23B0
`define TANH_LUT_POSITIVE_23B8 16'h23B8
`define TANH_LUT_POSITIVE_23C0 16'h23C0
`define TANH_LUT_POSITIVE_23C8 16'h23C8
`define TANH_LUT_POSITIVE_23D0 16'h23D0
`define TANH_LUT_POSITIVE_23D8 16'h23D8
`define TANH_LUT_POSITIVE_23E0 16'h23E0
`define TANH_LUT_POSITIVE_23E8 16'h23E8
`define TANH_LUT_POSITIVE_23F0 16'h23F0
`define TANH_LUT_POSITIVE_23F8 16'h23F8
`define TANH_LUT_POSITIVE_2400 16'h2400
`define TANH_LUT_POSITIVE_2408 16'h2408
`define TANH_LUT_POSITIVE_2410 16'h2410
`define TANH_LUT_POSITIVE_2418 16'h2418
`define TANH_LUT_POSITIVE_2420 16'h2420
`define TANH_LUT_POSITIVE_2428 16'h2428
`define TANH_LUT_POSITIVE_2430 16'h2430
`define TANH_LUT_POSITIVE_2438 16'h2438
`define TANH_LUT_POSITIVE_2440 16'h2440
`define TANH_LUT_POSITIVE_2448 16'h2448
`define TANH_LUT_POSITIVE_2450 16'h2450
`define TANH_LUT_POSITIVE_2458 16'h2458
`define TANH_LUT_POSITIVE_2460 16'h2460
`define TANH_LUT_POSITIVE_2468 16'h2468
`define TANH_LUT_POSITIVE_2470 16'h2470
`define TANH_LUT_POSITIVE_2478 16'h2478
`define TANH_LUT_POSITIVE_2480 16'h2480
`define TANH_LUT_POSITIVE_2488 16'h2488
`define TANH_LUT_POSITIVE_2490 16'h2490
`define TANH_LUT_POSITIVE_2498 16'h2498
`define TANH_LUT_POSITIVE_24A0 16'h24A0
`define TANH_LUT_POSITIVE_24A8 16'h24A8
`define TANH_LUT_POSITIVE_24B0 16'h24B0
`define TANH_LUT_POSITIVE_24B8 16'h24B8
`define TANH_LUT_POSITIVE_24C0 16'h24C0
`define TANH_LUT_POSITIVE_24C8 16'h24C8
`define TANH_LUT_POSITIVE_24D0 16'h24D0
`define TANH_LUT_POSITIVE_24D8 16'h24D8
`define TANH_LUT_POSITIVE_24E0 16'h24E0
`define TANH_LUT_POSITIVE_24E8 16'h24E8
`define TANH_LUT_POSITIVE_24F0 16'h24F0
`define TANH_LUT_POSITIVE_24F8 16'h24F8
`define TANH_LUT_POSITIVE_2500 16'h2500
`define TANH_LUT_POSITIVE_2508 16'h2508
`define TANH_LUT_POSITIVE_2510 16'h2510
`define TANH_LUT_POSITIVE_2518 16'h2518
`define TANH_LUT_POSITIVE_2520 16'h2520
`define TANH_LUT_POSITIVE_2528 16'h2528
`define TANH_LUT_POSITIVE_2530 16'h2530
`define TANH_LUT_POSITIVE_2538 16'h2538
`define TANH_LUT_POSITIVE_2540 16'h2540
`define TANH_LUT_POSITIVE_2548 16'h2548
`define TANH_LUT_POSITIVE_2550 16'h2550
`define TANH_LUT_POSITIVE_2558 16'h2558
`define TANH_LUT_POSITIVE_2560 16'h2560
`define TANH_LUT_POSITIVE_2568 16'h2568
`define TANH_LUT_POSITIVE_2570 16'h2570
`define TANH_LUT_POSITIVE_2578 16'h2578
`define TANH_LUT_POSITIVE_2580 16'h2580
`define TANH_LUT_POSITIVE_2588 16'h2588
`define TANH_LUT_POSITIVE_2590 16'h2590
`define TANH_LUT_POSITIVE_2598 16'h2598
`define TANH_LUT_POSITIVE_25A0 16'h25A0
`define TANH_LUT_POSITIVE_25A8 16'h25A8
`define TANH_LUT_POSITIVE_25B0 16'h25B0
`define TANH_LUT_POSITIVE_25B8 16'h25B8
`define TANH_LUT_POSITIVE_25C0 16'h25C0
`define TANH_LUT_POSITIVE_25C8 16'h25C8
`define TANH_LUT_POSITIVE_25D0 16'h25D0
`define TANH_LUT_POSITIVE_25D8 16'h25D8
`define TANH_LUT_POSITIVE_25E0 16'h25E0
`define TANH_LUT_POSITIVE_25E8 16'h25E8
`define TANH_LUT_POSITIVE_25F0 16'h25F0
`define TANH_LUT_POSITIVE_25F8 16'h25F8
`define TANH_LUT_POSITIVE_2600 16'h2600
`define TANH_LUT_POSITIVE_2608 16'h2608
`define TANH_LUT_POSITIVE_2610 16'h2610
`define TANH_LUT_POSITIVE_2618 16'h2618
`define TANH_LUT_POSITIVE_2620 16'h2620
`define TANH_LUT_POSITIVE_2628 16'h2628
`define TANH_LUT_POSITIVE_2630 16'h2630
`define TANH_LUT_POSITIVE_2638 16'h2638
`define TANH_LUT_POSITIVE_2640 16'h2640
`define TANH_LUT_POSITIVE_2648 16'h2648
`define TANH_LUT_POSITIVE_2650 16'h2650
`define TANH_LUT_POSITIVE_2658 16'h2658
`define TANH_LUT_POSITIVE_2660 16'h2660
`define TANH_LUT_POSITIVE_2668 16'h2668
`define TANH_LUT_POSITIVE_2670 16'h2670
`define TANH_LUT_POSITIVE_2678 16'h2678
`define TANH_LUT_POSITIVE_2680 16'h2680
`define TANH_LUT_POSITIVE_2688 16'h2688
`define TANH_LUT_POSITIVE_2690 16'h2690
`define TANH_LUT_POSITIVE_2698 16'h2698
`define TANH_LUT_POSITIVE_26A0 16'h26A0
`define TANH_LUT_POSITIVE_26A8 16'h26A8
`define TANH_LUT_POSITIVE_26B0 16'h26B0
`define TANH_LUT_POSITIVE_26B8 16'h26B8
`define TANH_LUT_POSITIVE_26C0 16'h26C0
`define TANH_LUT_POSITIVE_26C8 16'h26C8
`define TANH_LUT_POSITIVE_26D0 16'h26D0
`define TANH_LUT_POSITIVE_26D8 16'h26D8
`define TANH_LUT_POSITIVE_26E0 16'h26E0
`define TANH_LUT_POSITIVE_26E8 16'h26E8
`define TANH_LUT_POSITIVE_26F0 16'h26F0
`define TANH_LUT_POSITIVE_26F8 16'h26F8
`define TANH_LUT_POSITIVE_2700 16'h2700
`define TANH_LUT_POSITIVE_2708 16'h2708
`define TANH_LUT_POSITIVE_2710 16'h2710
`define TANH_LUT_POSITIVE_2718 16'h2718
`define TANH_LUT_POSITIVE_2720 16'h2720
`define TANH_LUT_POSITIVE_2728 16'h2728
`define TANH_LUT_POSITIVE_2730 16'h2730
`define TANH_LUT_POSITIVE_2738 16'h2738
`define TANH_LUT_POSITIVE_2740 16'h2740
`define TANH_LUT_POSITIVE_2748 16'h2747
`define TANH_LUT_POSITIVE_2750 16'h274F
`define TANH_LUT_POSITIVE_2758 16'h2757
`define TANH_LUT_POSITIVE_2760 16'h275F
`define TANH_LUT_POSITIVE_2768 16'h2767
`define TANH_LUT_POSITIVE_2770 16'h276F
`define TANH_LUT_POSITIVE_2778 16'h2777
`define TANH_LUT_POSITIVE_2780 16'h277F
`define TANH_LUT_POSITIVE_2788 16'h2787
`define TANH_LUT_POSITIVE_2790 16'h278F
`define TANH_LUT_POSITIVE_2798 16'h2797
`define TANH_LUT_POSITIVE_27A0 16'h279F
`define TANH_LUT_POSITIVE_27A8 16'h27A7
`define TANH_LUT_POSITIVE_27B0 16'h27AF
`define TANH_LUT_POSITIVE_27B8 16'h27B7
`define TANH_LUT_POSITIVE_27C0 16'h27BF
`define TANH_LUT_POSITIVE_27C8 16'h27C7
`define TANH_LUT_POSITIVE_27D0 16'h27CF
`define TANH_LUT_POSITIVE_27D8 16'h27D7
`define TANH_LUT_POSITIVE_27E0 16'h27DF
`define TANH_LUT_POSITIVE_27E8 16'h27E7
`define TANH_LUT_POSITIVE_27F0 16'h27EF
`define TANH_LUT_POSITIVE_27F8 16'h27F7
`define TANH_LUT_POSITIVE_2800 16'h27FF
`define TANH_LUT_POSITIVE_2808 16'h2808
`define TANH_LUT_POSITIVE_2810 16'h2810
`define TANH_LUT_POSITIVE_2818 16'h2818
`define TANH_LUT_POSITIVE_2820 16'h2820
`define TANH_LUT_POSITIVE_2828 16'h2828
`define TANH_LUT_POSITIVE_2830 16'h2830
`define TANH_LUT_POSITIVE_2838 16'h2838
`define TANH_LUT_POSITIVE_2840 16'h2840
`define TANH_LUT_POSITIVE_2848 16'h2848
`define TANH_LUT_POSITIVE_2850 16'h2850
`define TANH_LUT_POSITIVE_2858 16'h2858
`define TANH_LUT_POSITIVE_2860 16'h2860
`define TANH_LUT_POSITIVE_2868 16'h2868
`define TANH_LUT_POSITIVE_2870 16'h2870
`define TANH_LUT_POSITIVE_2878 16'h2878
`define TANH_LUT_POSITIVE_2880 16'h2880
`define TANH_LUT_POSITIVE_2888 16'h2888
`define TANH_LUT_POSITIVE_2890 16'h2890
`define TANH_LUT_POSITIVE_2898 16'h2897
`define TANH_LUT_POSITIVE_28A0 16'h289F
`define TANH_LUT_POSITIVE_28A8 16'h28A7
`define TANH_LUT_POSITIVE_28B0 16'h28AF
`define TANH_LUT_POSITIVE_28B8 16'h28B7
`define TANH_LUT_POSITIVE_28C0 16'h28BF
`define TANH_LUT_POSITIVE_28C8 16'h28C7
`define TANH_LUT_POSITIVE_28D0 16'h28CF
`define TANH_LUT_POSITIVE_28D8 16'h28D7
`define TANH_LUT_POSITIVE_28E0 16'h28DF
`define TANH_LUT_POSITIVE_28E8 16'h28E7
`define TANH_LUT_POSITIVE_28F0 16'h28EF
`define TANH_LUT_POSITIVE_28F8 16'h28F7
`define TANH_LUT_POSITIVE_2900 16'h28FF
`define TANH_LUT_POSITIVE_2908 16'h2907
`define TANH_LUT_POSITIVE_2910 16'h290F
`define TANH_LUT_POSITIVE_2918 16'h2917
`define TANH_LUT_POSITIVE_2920 16'h291F
`define TANH_LUT_POSITIVE_2928 16'h2927
`define TANH_LUT_POSITIVE_2930 16'h292F
`define TANH_LUT_POSITIVE_2938 16'h2937
`define TANH_LUT_POSITIVE_2940 16'h293F
`define TANH_LUT_POSITIVE_2948 16'h2947
`define TANH_LUT_POSITIVE_2950 16'h294F
`define TANH_LUT_POSITIVE_2958 16'h2957
`define TANH_LUT_POSITIVE_2960 16'h295F
`define TANH_LUT_POSITIVE_2968 16'h2967
`define TANH_LUT_POSITIVE_2970 16'h296F
`define TANH_LUT_POSITIVE_2978 16'h2977
`define TANH_LUT_POSITIVE_2980 16'h297F
`define TANH_LUT_POSITIVE_2988 16'h2987
`define TANH_LUT_POSITIVE_2990 16'h298F
`define TANH_LUT_POSITIVE_2998 16'h2997
`define TANH_LUT_POSITIVE_29A0 16'h299F
`define TANH_LUT_POSITIVE_29A8 16'h29A7
`define TANH_LUT_POSITIVE_29B0 16'h29AF
`define TANH_LUT_POSITIVE_29B8 16'h29B7
`define TANH_LUT_POSITIVE_29C0 16'h29BF
`define TANH_LUT_POSITIVE_29C8 16'h29C7
`define TANH_LUT_POSITIVE_29D0 16'h29CF
`define TANH_LUT_POSITIVE_29D8 16'h29D7
`define TANH_LUT_POSITIVE_29E0 16'h29DF
`define TANH_LUT_POSITIVE_29E8 16'h29E7
`define TANH_LUT_POSITIVE_29F0 16'h29EF
`define TANH_LUT_POSITIVE_29F8 16'h29F7
`define TANH_LUT_POSITIVE_2A00 16'h29FF
`define TANH_LUT_POSITIVE_2A08 16'h2A07
`define TANH_LUT_POSITIVE_2A10 16'h2A0F
`define TANH_LUT_POSITIVE_2A18 16'h2A17
`define TANH_LUT_POSITIVE_2A20 16'h2A1F
`define TANH_LUT_POSITIVE_2A28 16'h2A27
`define TANH_LUT_POSITIVE_2A30 16'h2A2F
`define TANH_LUT_POSITIVE_2A38 16'h2A37
`define TANH_LUT_POSITIVE_2A40 16'h2A3F
`define TANH_LUT_POSITIVE_2A48 16'h2A47
`define TANH_LUT_POSITIVE_2A50 16'h2A4F
`define TANH_LUT_POSITIVE_2A58 16'h2A57
`define TANH_LUT_POSITIVE_2A60 16'h2A5F
`define TANH_LUT_POSITIVE_2A68 16'h2A67
`define TANH_LUT_POSITIVE_2A70 16'h2A6F
`define TANH_LUT_POSITIVE_2A78 16'h2A77
`define TANH_LUT_POSITIVE_2A80 16'h2A7F
`define TANH_LUT_POSITIVE_2A88 16'h2A87
`define TANH_LUT_POSITIVE_2A90 16'h2A8F
`define TANH_LUT_POSITIVE_2A98 16'h2A97
`define TANH_LUT_POSITIVE_2AA0 16'h2A9E
`define TANH_LUT_POSITIVE_2AA8 16'h2AA6
`define TANH_LUT_POSITIVE_2AB0 16'h2AAE
`define TANH_LUT_POSITIVE_2AB8 16'h2AB6
`define TANH_LUT_POSITIVE_2AC0 16'h2ABE
`define TANH_LUT_POSITIVE_2AC8 16'h2AC6
`define TANH_LUT_POSITIVE_2AD0 16'h2ACE
`define TANH_LUT_POSITIVE_2AD8 16'h2AD6
`define TANH_LUT_POSITIVE_2AE0 16'h2ADE
`define TANH_LUT_POSITIVE_2AE8 16'h2AE6
`define TANH_LUT_POSITIVE_2AF0 16'h2AEE
`define TANH_LUT_POSITIVE_2AF8 16'h2AF6
`define TANH_LUT_POSITIVE_2B00 16'h2AFE
`define TANH_LUT_POSITIVE_2B08 16'h2B06
`define TANH_LUT_POSITIVE_2B10 16'h2B0E
`define TANH_LUT_POSITIVE_2B18 16'h2B16
`define TANH_LUT_POSITIVE_2B20 16'h2B1E
`define TANH_LUT_POSITIVE_2B28 16'h2B26
`define TANH_LUT_POSITIVE_2B30 16'h2B2E
`define TANH_LUT_POSITIVE_2B38 16'h2B36
`define TANH_LUT_POSITIVE_2B40 16'h2B3E
`define TANH_LUT_POSITIVE_2B48 16'h2B46
`define TANH_LUT_POSITIVE_2B50 16'h2B4E
`define TANH_LUT_POSITIVE_2B58 16'h2B56
`define TANH_LUT_POSITIVE_2B60 16'h2B5E
`define TANH_LUT_POSITIVE_2B68 16'h2B66
`define TANH_LUT_POSITIVE_2B70 16'h2B6E
`define TANH_LUT_POSITIVE_2B78 16'h2B76
`define TANH_LUT_POSITIVE_2B80 16'h2B7E
`define TANH_LUT_POSITIVE_2B88 16'h2B86
`define TANH_LUT_POSITIVE_2B90 16'h2B8E
`define TANH_LUT_POSITIVE_2B98 16'h2B96
`define TANH_LUT_POSITIVE_2BA0 16'h2B9E
`define TANH_LUT_POSITIVE_2BA8 16'h2BA6
`define TANH_LUT_POSITIVE_2BB0 16'h2BAE
`define TANH_LUT_POSITIVE_2BB8 16'h2BB6
`define TANH_LUT_POSITIVE_2BC0 16'h2BBE
`define TANH_LUT_POSITIVE_2BC8 16'h2BC6
`define TANH_LUT_POSITIVE_2BD0 16'h2BCE
`define TANH_LUT_POSITIVE_2BD8 16'h2BD5
`define TANH_LUT_POSITIVE_2BE0 16'h2BDD
`define TANH_LUT_POSITIVE_2BE8 16'h2BE5
`define TANH_LUT_POSITIVE_2BF0 16'h2BED
`define TANH_LUT_POSITIVE_2BF8 16'h2BF5
`define TANH_LUT_POSITIVE_2C00 16'h2BFD
`define TANH_LUT_POSITIVE_2C08 16'h2C07
`define TANH_LUT_POSITIVE_2C10 16'h2C0F
`define TANH_LUT_POSITIVE_2C18 16'h2C17
`define TANH_LUT_POSITIVE_2C20 16'h2C1F
`define TANH_LUT_POSITIVE_2C28 16'h2C27
`define TANH_LUT_POSITIVE_2C30 16'h2C2E
`define TANH_LUT_POSITIVE_2C38 16'h2C36
`define TANH_LUT_POSITIVE_2C40 16'h2C3E
`define TANH_LUT_POSITIVE_2C48 16'h2C46
`define TANH_LUT_POSITIVE_2C50 16'h2C4E
`define TANH_LUT_POSITIVE_2C58 16'h2C56
`define TANH_LUT_POSITIVE_2C60 16'h2C5E
`define TANH_LUT_POSITIVE_2C68 16'h2C66
`define TANH_LUT_POSITIVE_2C70 16'h2C6E
`define TANH_LUT_POSITIVE_2C78 16'h2C76
`define TANH_LUT_POSITIVE_2C80 16'h2C7E
`define TANH_LUT_POSITIVE_2C88 16'h2C86
`define TANH_LUT_POSITIVE_2C90 16'h2C8E
`define TANH_LUT_POSITIVE_2C98 16'h2C96
`define TANH_LUT_POSITIVE_2CA0 16'h2C9E
`define TANH_LUT_POSITIVE_2CA8 16'h2CA6
`define TANH_LUT_POSITIVE_2CB0 16'h2CAE
`define TANH_LUT_POSITIVE_2CB8 16'h2CB6
`define TANH_LUT_POSITIVE_2CC0 16'h2CBE
`define TANH_LUT_POSITIVE_2CC8 16'h2CC6
`define TANH_LUT_POSITIVE_2CD0 16'h2CCE
`define TANH_LUT_POSITIVE_2CD8 16'h2CD6
`define TANH_LUT_POSITIVE_2CE0 16'h2CDE
`define TANH_LUT_POSITIVE_2CE8 16'h2CE6
`define TANH_LUT_POSITIVE_2CF0 16'h2CED
`define TANH_LUT_POSITIVE_2CF8 16'h2CF5
`define TANH_LUT_POSITIVE_2D00 16'h2CFD
`define TANH_LUT_POSITIVE_2D08 16'h2D05
`define TANH_LUT_POSITIVE_2D10 16'h2D0D
`define TANH_LUT_POSITIVE_2D18 16'h2D15
`define TANH_LUT_POSITIVE_2D20 16'h2D1D
`define TANH_LUT_POSITIVE_2D28 16'h2D25
`define TANH_LUT_POSITIVE_2D30 16'h2D2D
`define TANH_LUT_POSITIVE_2D38 16'h2D35
`define TANH_LUT_POSITIVE_2D40 16'h2D3D
`define TANH_LUT_POSITIVE_2D48 16'h2D45
`define TANH_LUT_POSITIVE_2D50 16'h2D4D
`define TANH_LUT_POSITIVE_2D58 16'h2D55
`define TANH_LUT_POSITIVE_2D60 16'h2D5D
`define TANH_LUT_POSITIVE_2D68 16'h2D65
`define TANH_LUT_POSITIVE_2D70 16'h2D6D
`define TANH_LUT_POSITIVE_2D78 16'h2D75
`define TANH_LUT_POSITIVE_2D80 16'h2D7D
`define TANH_LUT_POSITIVE_2D88 16'h2D84
`define TANH_LUT_POSITIVE_2D90 16'h2D8C
`define TANH_LUT_POSITIVE_2D98 16'h2D94
`define TANH_LUT_POSITIVE_2DA0 16'h2D9C
`define TANH_LUT_POSITIVE_2DA8 16'h2DA4
`define TANH_LUT_POSITIVE_2DB0 16'h2DAC
`define TANH_LUT_POSITIVE_2DB8 16'h2DB4
`define TANH_LUT_POSITIVE_2DC0 16'h2DBC
`define TANH_LUT_POSITIVE_2DC8 16'h2DC4
`define TANH_LUT_POSITIVE_2DD0 16'h2DCC
`define TANH_LUT_POSITIVE_2DD8 16'h2DD4
`define TANH_LUT_POSITIVE_2DE0 16'h2DDC
`define TANH_LUT_POSITIVE_2DE8 16'h2DE4
`define TANH_LUT_POSITIVE_2DF0 16'h2DEC
`define TANH_LUT_POSITIVE_2DF8 16'h2DF4
`define TANH_LUT_POSITIVE_2E00 16'h2DFC
`define TANH_LUT_POSITIVE_2E08 16'h2E03
`define TANH_LUT_POSITIVE_2E10 16'h2E0B
`define TANH_LUT_POSITIVE_2E18 16'h2E13
`define TANH_LUT_POSITIVE_2E20 16'h2E1B
`define TANH_LUT_POSITIVE_2E28 16'h2E23
`define TANH_LUT_POSITIVE_2E30 16'h2E2B
`define TANH_LUT_POSITIVE_2E38 16'h2E33
`define TANH_LUT_POSITIVE_2E40 16'h2E3B
`define TANH_LUT_POSITIVE_2E48 16'h2E43
`define TANH_LUT_POSITIVE_2E50 16'h2E4B
`define TANH_LUT_POSITIVE_2E58 16'h2E53
`define TANH_LUT_POSITIVE_2E60 16'h2E5B
`define TANH_LUT_POSITIVE_2E68 16'h2E63
`define TANH_LUT_POSITIVE_2E70 16'h2E6A
`define TANH_LUT_POSITIVE_2E78 16'h2E72
`define TANH_LUT_POSITIVE_2E80 16'h2E7A
`define TANH_LUT_POSITIVE_2E88 16'h2E82
`define TANH_LUT_POSITIVE_2E90 16'h2E8A
`define TANH_LUT_POSITIVE_2E98 16'h2E92
`define TANH_LUT_POSITIVE_2EA0 16'h2E9A
`define TANH_LUT_POSITIVE_2EA8 16'h2EA2
`define TANH_LUT_POSITIVE_2EB0 16'h2EAA
`define TANH_LUT_POSITIVE_2EB8 16'h2EB2
`define TANH_LUT_POSITIVE_2EC0 16'h2EBA
`define TANH_LUT_POSITIVE_2EC8 16'h2EC2
`define TANH_LUT_POSITIVE_2ED0 16'h2EC9
`define TANH_LUT_POSITIVE_2ED8 16'h2ED1
`define TANH_LUT_POSITIVE_2EE0 16'h2ED9
`define TANH_LUT_POSITIVE_2EE8 16'h2EE1
`define TANH_LUT_POSITIVE_2EF0 16'h2EE9
`define TANH_LUT_POSITIVE_2EF8 16'h2EF1
`define TANH_LUT_POSITIVE_2F00 16'h2EF9
`define TANH_LUT_POSITIVE_2F08 16'h2F01
`define TANH_LUT_POSITIVE_2F10 16'h2F09
`define TANH_LUT_POSITIVE_2F18 16'h2F11
`define TANH_LUT_POSITIVE_2F20 16'h2F19
`define TANH_LUT_POSITIVE_2F28 16'h2F20
`define TANH_LUT_POSITIVE_2F30 16'h2F28
`define TANH_LUT_POSITIVE_2F38 16'h2F30
`define TANH_LUT_POSITIVE_2F40 16'h2F38
`define TANH_LUT_POSITIVE_2F48 16'h2F40
`define TANH_LUT_POSITIVE_2F50 16'h2F48
`define TANH_LUT_POSITIVE_2F58 16'h2F50
`define TANH_LUT_POSITIVE_2F60 16'h2F58
`define TANH_LUT_POSITIVE_2F68 16'h2F60
`define TANH_LUT_POSITIVE_2F70 16'h2F67
`define TANH_LUT_POSITIVE_2F78 16'h2F6F
`define TANH_LUT_POSITIVE_2F80 16'h2F77
`define TANH_LUT_POSITIVE_2F88 16'h2F7F
`define TANH_LUT_POSITIVE_2F90 16'h2F87
`define TANH_LUT_POSITIVE_2F98 16'h2F8F
`define TANH_LUT_POSITIVE_2FA0 16'h2F97
`define TANH_LUT_POSITIVE_2FA8 16'h2F9F
`define TANH_LUT_POSITIVE_2FB0 16'h2FA7
`define TANH_LUT_POSITIVE_2FB8 16'h2FAE
`define TANH_LUT_POSITIVE_2FC0 16'h2FB6
`define TANH_LUT_POSITIVE_2FC8 16'h2FBE
`define TANH_LUT_POSITIVE_2FD0 16'h2FC6
`define TANH_LUT_POSITIVE_2FD8 16'h2FCE
`define TANH_LUT_POSITIVE_2FE0 16'h2FD6
`define TANH_LUT_POSITIVE_2FE8 16'h2FDE
`define TANH_LUT_POSITIVE_2FF0 16'h2FE6
`define TANH_LUT_POSITIVE_2FF8 16'h2FEE
`define TANH_LUT_POSITIVE_3000 16'h2FF5
`define TANH_LUT_POSITIVE_3008 16'h3003
`define TANH_LUT_POSITIVE_3010 16'h300A
`define TANH_LUT_POSITIVE_3018 16'h3012
`define TANH_LUT_POSITIVE_3020 16'h301A
`define TANH_LUT_POSITIVE_3028 16'h3022
`define TANH_LUT_POSITIVE_3030 16'h302A
`define TANH_LUT_POSITIVE_3038 16'h3032
`define TANH_LUT_POSITIVE_3040 16'h303A
`define TANH_LUT_POSITIVE_3048 16'h3042
`define TANH_LUT_POSITIVE_3050 16'h3049
`define TANH_LUT_POSITIVE_3058 16'h3051
`define TANH_LUT_POSITIVE_3060 16'h3059
`define TANH_LUT_POSITIVE_3068 16'h3061
`define TANH_LUT_POSITIVE_3070 16'h3069
`define TANH_LUT_POSITIVE_3078 16'h3071
`define TANH_LUT_POSITIVE_3080 16'h3078
`define TANH_LUT_POSITIVE_3088 16'h3080
`define TANH_LUT_POSITIVE_3090 16'h3088
`define TANH_LUT_POSITIVE_3098 16'h3090
`define TANH_LUT_POSITIVE_30A0 16'h3098
`define TANH_LUT_POSITIVE_30A8 16'h30A0
`define TANH_LUT_POSITIVE_30B0 16'h30A7
`define TANH_LUT_POSITIVE_30B8 16'h30AF
`define TANH_LUT_POSITIVE_30C0 16'h30B7
`define TANH_LUT_POSITIVE_30C8 16'h30BF
`define TANH_LUT_POSITIVE_30D0 16'h30C7
`define TANH_LUT_POSITIVE_30D8 16'h30CF
`define TANH_LUT_POSITIVE_30E0 16'h30D6
`define TANH_LUT_POSITIVE_30E8 16'h30DE
`define TANH_LUT_POSITIVE_30F0 16'h30E6
`define TANH_LUT_POSITIVE_30F8 16'h30EE
`define TANH_LUT_POSITIVE_3100 16'h30F6
`define TANH_LUT_POSITIVE_3108 16'h30FD
`define TANH_LUT_POSITIVE_3110 16'h3105
`define TANH_LUT_POSITIVE_3118 16'h310D
`define TANH_LUT_POSITIVE_3120 16'h3115
`define TANH_LUT_POSITIVE_3128 16'h311D
`define TANH_LUT_POSITIVE_3130 16'h3124
`define TANH_LUT_POSITIVE_3138 16'h312C
`define TANH_LUT_POSITIVE_3140 16'h3134
`define TANH_LUT_POSITIVE_3148 16'h313C
`define TANH_LUT_POSITIVE_3150 16'h3144
`define TANH_LUT_POSITIVE_3158 16'h314B
`define TANH_LUT_POSITIVE_3160 16'h3153
`define TANH_LUT_POSITIVE_3168 16'h315B
`define TANH_LUT_POSITIVE_3170 16'h3163
`define TANH_LUT_POSITIVE_3178 16'h316B
`define TANH_LUT_POSITIVE_3180 16'h3172
`define TANH_LUT_POSITIVE_3188 16'h317A
`define TANH_LUT_POSITIVE_3190 16'h3182
`define TANH_LUT_POSITIVE_3198 16'h318A
`define TANH_LUT_POSITIVE_31A0 16'h3191
`define TANH_LUT_POSITIVE_31A8 16'h3199
`define TANH_LUT_POSITIVE_31B0 16'h31A1
`define TANH_LUT_POSITIVE_31B8 16'h31A9
`define TANH_LUT_POSITIVE_31C0 16'h31B0
`define TANH_LUT_POSITIVE_31C8 16'h31B8
`define TANH_LUT_POSITIVE_31D0 16'h31C0
`define TANH_LUT_POSITIVE_31D8 16'h31C8
`define TANH_LUT_POSITIVE_31E0 16'h31CF
`define TANH_LUT_POSITIVE_31E8 16'h31D7
`define TANH_LUT_POSITIVE_31F0 16'h31DF
`define TANH_LUT_POSITIVE_31F8 16'h31E7
`define TANH_LUT_POSITIVE_3200 16'h31EE
`define TANH_LUT_POSITIVE_3208 16'h31F6
`define TANH_LUT_POSITIVE_3210 16'h31FE
`define TANH_LUT_POSITIVE_3218 16'h3205
`define TANH_LUT_POSITIVE_3220 16'h320D
`define TANH_LUT_POSITIVE_3228 16'h3215
`define TANH_LUT_POSITIVE_3230 16'h321D
`define TANH_LUT_POSITIVE_3238 16'h3224
`define TANH_LUT_POSITIVE_3240 16'h322C
`define TANH_LUT_POSITIVE_3248 16'h3234
`define TANH_LUT_POSITIVE_3250 16'h323B
`define TANH_LUT_POSITIVE_3258 16'h3243
`define TANH_LUT_POSITIVE_3260 16'h324B
`define TANH_LUT_POSITIVE_3268 16'h3252
`define TANH_LUT_POSITIVE_3270 16'h325A
`define TANH_LUT_POSITIVE_3278 16'h3262
`define TANH_LUT_POSITIVE_3280 16'h3269
`define TANH_LUT_POSITIVE_3288 16'h3271
`define TANH_LUT_POSITIVE_3290 16'h3279
`define TANH_LUT_POSITIVE_3298 16'h3281
`define TANH_LUT_POSITIVE_32A0 16'h3288
`define TANH_LUT_POSITIVE_32A8 16'h3290
`define TANH_LUT_POSITIVE_32B0 16'h3298
`define TANH_LUT_POSITIVE_32B8 16'h329F
`define TANH_LUT_POSITIVE_32C0 16'h32A7
`define TANH_LUT_POSITIVE_32C8 16'h32AE
`define TANH_LUT_POSITIVE_32D0 16'h32B6
`define TANH_LUT_POSITIVE_32D8 16'h32BE
`define TANH_LUT_POSITIVE_32E0 16'h32C5
`define TANH_LUT_POSITIVE_32E8 16'h32CD
`define TANH_LUT_POSITIVE_32F0 16'h32D5
`define TANH_LUT_POSITIVE_32F8 16'h32DC
`define TANH_LUT_POSITIVE_3300 16'h32E4
`define TANH_LUT_POSITIVE_3308 16'h32EC
`define TANH_LUT_POSITIVE_3310 16'h32F3
`define TANH_LUT_POSITIVE_3318 16'h32FB
`define TANH_LUT_POSITIVE_3320 16'h3302
`define TANH_LUT_POSITIVE_3328 16'h330A
`define TANH_LUT_POSITIVE_3330 16'h3312
`define TANH_LUT_POSITIVE_3338 16'h3319
`define TANH_LUT_POSITIVE_3340 16'h3321
`define TANH_LUT_POSITIVE_3348 16'h3328
`define TANH_LUT_POSITIVE_3350 16'h3330
`define TANH_LUT_POSITIVE_3358 16'h3338
`define TANH_LUT_POSITIVE_3360 16'h333F
`define TANH_LUT_POSITIVE_3368 16'h3347
`define TANH_LUT_POSITIVE_3370 16'h334E
`define TANH_LUT_POSITIVE_3378 16'h3356
`define TANH_LUT_POSITIVE_3380 16'h335E
`define TANH_LUT_POSITIVE_3388 16'h3365
`define TANH_LUT_POSITIVE_3390 16'h336D
`define TANH_LUT_POSITIVE_3398 16'h3374
`define TANH_LUT_POSITIVE_33A0 16'h337C
`define TANH_LUT_POSITIVE_33A8 16'h3383
`define TANH_LUT_POSITIVE_33B0 16'h338B
`define TANH_LUT_POSITIVE_33B8 16'h3393
`define TANH_LUT_POSITIVE_33C0 16'h339A
`define TANH_LUT_POSITIVE_33C8 16'h33A2
`define TANH_LUT_POSITIVE_33D0 16'h33A9
`define TANH_LUT_POSITIVE_33D8 16'h33B1
`define TANH_LUT_POSITIVE_33E0 16'h33B8
`define TANH_LUT_POSITIVE_33E8 16'h33C0
`define TANH_LUT_POSITIVE_33F0 16'h33C7
`define TANH_LUT_POSITIVE_33F8 16'h33CF
`define TANH_LUT_POSITIVE_3400 16'h33D6
`define TANH_LUT_POSITIVE_3408 16'h33E5
`define TANH_LUT_POSITIVE_3410 16'h33F4
`define TANH_LUT_POSITIVE_3418 16'h3402
`define TANH_LUT_POSITIVE_3420 16'h3409
`define TANH_LUT_POSITIVE_3428 16'h3411
`define TANH_LUT_POSITIVE_3430 16'h3418
`define TANH_LUT_POSITIVE_3438 16'h3420
`define TANH_LUT_POSITIVE_3440 16'h3427
`define TANH_LUT_POSITIVE_3448 16'h342F
`define TANH_LUT_POSITIVE_3450 16'h3436
`define TANH_LUT_POSITIVE_3458 16'h343D
`define TANH_LUT_POSITIVE_3460 16'h3445
`define TANH_LUT_POSITIVE_3468 16'h344C
`define TANH_LUT_POSITIVE_3470 16'h3454
`define TANH_LUT_POSITIVE_3478 16'h345B
`define TANH_LUT_POSITIVE_3480 16'h3463
`define TANH_LUT_POSITIVE_3488 16'h346A
`define TANH_LUT_POSITIVE_3490 16'h3471
`define TANH_LUT_POSITIVE_3498 16'h3479
`define TANH_LUT_POSITIVE_34A0 16'h3480
`define TANH_LUT_POSITIVE_34A8 16'h3487
`define TANH_LUT_POSITIVE_34B0 16'h348F
`define TANH_LUT_POSITIVE_34B8 16'h3496
`define TANH_LUT_POSITIVE_34C0 16'h349D
`define TANH_LUT_POSITIVE_34C8 16'h34A5
`define TANH_LUT_POSITIVE_34D0 16'h34AC
`define TANH_LUT_POSITIVE_34D8 16'h34B3
`define TANH_LUT_POSITIVE_34E0 16'h34BB
`define TANH_LUT_POSITIVE_34E8 16'h34C2
`define TANH_LUT_POSITIVE_34F0 16'h34C9
`define TANH_LUT_POSITIVE_34F8 16'h34D1
`define TANH_LUT_POSITIVE_3500 16'h34D8
`define TANH_LUT_POSITIVE_3508 16'h34DF
`define TANH_LUT_POSITIVE_3510 16'h34E6
`define TANH_LUT_POSITIVE_3518 16'h34EE
`define TANH_LUT_POSITIVE_3520 16'h34F5
`define TANH_LUT_POSITIVE_3528 16'h34FC
`define TANH_LUT_POSITIVE_3530 16'h3503
`define TANH_LUT_POSITIVE_3538 16'h350B
`define TANH_LUT_POSITIVE_3540 16'h3512
`define TANH_LUT_POSITIVE_3548 16'h3519
`define TANH_LUT_POSITIVE_3550 16'h3520
`define TANH_LUT_POSITIVE_3558 16'h3527
`define TANH_LUT_POSITIVE_3560 16'h352E
`define TANH_LUT_POSITIVE_3568 16'h3536
`define TANH_LUT_POSITIVE_3570 16'h353D
`define TANH_LUT_POSITIVE_3578 16'h3544
`define TANH_LUT_POSITIVE_3580 16'h354B
`define TANH_LUT_POSITIVE_3588 16'h3552
`define TANH_LUT_POSITIVE_3590 16'h3559
`define TANH_LUT_POSITIVE_3598 16'h3560
`define TANH_LUT_POSITIVE_35A0 16'h3567
`define TANH_LUT_POSITIVE_35A8 16'h356F
`define TANH_LUT_POSITIVE_35B0 16'h3576
`define TANH_LUT_POSITIVE_35B8 16'h357D
`define TANH_LUT_POSITIVE_35C0 16'h3584
`define TANH_LUT_POSITIVE_35C8 16'h358B
`define TANH_LUT_POSITIVE_35D0 16'h3592
`define TANH_LUT_POSITIVE_35D8 16'h3599
`define TANH_LUT_POSITIVE_35E0 16'h35A0
`define TANH_LUT_POSITIVE_35E8 16'h35A7
`define TANH_LUT_POSITIVE_35F0 16'h35AE
`define TANH_LUT_POSITIVE_35F8 16'h35B5
`define TANH_LUT_POSITIVE_3600 16'h35BC
`define TANH_LUT_POSITIVE_3608 16'h35C3
`define TANH_LUT_POSITIVE_3610 16'h35CA
`define TANH_LUT_POSITIVE_3618 16'h35D1
`define TANH_LUT_POSITIVE_3620 16'h35D8
`define TANH_LUT_POSITIVE_3628 16'h35DF
`define TANH_LUT_POSITIVE_3630 16'h35E5
`define TANH_LUT_POSITIVE_3638 16'h35EC
`define TANH_LUT_POSITIVE_3640 16'h35F3
`define TANH_LUT_POSITIVE_3648 16'h35FA
`define TANH_LUT_POSITIVE_3650 16'h3601
`define TANH_LUT_POSITIVE_3658 16'h3608
`define TANH_LUT_POSITIVE_3660 16'h360F
`define TANH_LUT_POSITIVE_3668 16'h3616
`define TANH_LUT_POSITIVE_3670 16'h361C
`define TANH_LUT_POSITIVE_3678 16'h3623
`define TANH_LUT_POSITIVE_3680 16'h362A
`define TANH_LUT_POSITIVE_3688 16'h3631
`define TANH_LUT_POSITIVE_3690 16'h3638
`define TANH_LUT_POSITIVE_3698 16'h363F
`define TANH_LUT_POSITIVE_36A0 16'h3645
`define TANH_LUT_POSITIVE_36A8 16'h364C
`define TANH_LUT_POSITIVE_36B0 16'h3653
`define TANH_LUT_POSITIVE_36B8 16'h365A
`define TANH_LUT_POSITIVE_36C0 16'h3660
`define TANH_LUT_POSITIVE_36C8 16'h3667
`define TANH_LUT_POSITIVE_36D0 16'h366E
`define TANH_LUT_POSITIVE_36D8 16'h3674
`define TANH_LUT_POSITIVE_36E0 16'h367B
`define TANH_LUT_POSITIVE_36E8 16'h3682
`define TANH_LUT_POSITIVE_36F0 16'h3688
`define TANH_LUT_POSITIVE_36F8 16'h368F
`define TANH_LUT_POSITIVE_3700 16'h3696
`define TANH_LUT_POSITIVE_3708 16'h369C
`define TANH_LUT_POSITIVE_3710 16'h36A3
`define TANH_LUT_POSITIVE_3718 16'h36AA
`define TANH_LUT_POSITIVE_3720 16'h36B0
`define TANH_LUT_POSITIVE_3728 16'h36B7
`define TANH_LUT_POSITIVE_3730 16'h36BD
`define TANH_LUT_POSITIVE_3738 16'h36C4
`define TANH_LUT_POSITIVE_3740 16'h36CB
`define TANH_LUT_POSITIVE_3748 16'h36D1
`define TANH_LUT_POSITIVE_3750 16'h36D8
`define TANH_LUT_POSITIVE_3758 16'h36DE
`define TANH_LUT_POSITIVE_3760 16'h36E5
`define TANH_LUT_POSITIVE_3768 16'h36EB
`define TANH_LUT_POSITIVE_3770 16'h36F2
`define TANH_LUT_POSITIVE_3778 16'h36F8
`define TANH_LUT_POSITIVE_3780 16'h36FF
`define TANH_LUT_POSITIVE_3788 16'h3705
`define TANH_LUT_POSITIVE_3790 16'h370C
`define TANH_LUT_POSITIVE_3798 16'h3712
`define TANH_LUT_POSITIVE_37A0 16'h3719
`define TANH_LUT_POSITIVE_37A8 16'h371F
`define TANH_LUT_POSITIVE_37B0 16'h3725
`define TANH_LUT_POSITIVE_37B8 16'h372C
`define TANH_LUT_POSITIVE_37C0 16'h3732
`define TANH_LUT_POSITIVE_37C8 16'h3739
`define TANH_LUT_POSITIVE_37D0 16'h373F
`define TANH_LUT_POSITIVE_37D8 16'h3745
`define TANH_LUT_POSITIVE_37E0 16'h374C
`define TANH_LUT_POSITIVE_37E8 16'h3752
`define TANH_LUT_POSITIVE_37F0 16'h3758
`define TANH_LUT_POSITIVE_37F8 16'h375F
`define TANH_LUT_POSITIVE_3800 16'h3765
`define TANH_LUT_POSITIVE_3808 16'h3771
`define TANH_LUT_POSITIVE_3810 16'h377E
`define TANH_LUT_POSITIVE_3818 16'h378A
`define TANH_LUT_POSITIVE_3820 16'h3797
`define TANH_LUT_POSITIVE_3828 16'h37A3
`define TANH_LUT_POSITIVE_3830 16'h37B0
`define TANH_LUT_POSITIVE_3838 16'h37BC
`define TANH_LUT_POSITIVE_3840 16'h37C8
`define TANH_LUT_POSITIVE_3848 16'h37D4
`define TANH_LUT_POSITIVE_3850 16'h37E0
`define TANH_LUT_POSITIVE_3858 16'h37EC
`define TANH_LUT_POSITIVE_3860 16'h37F9
`define TANH_LUT_POSITIVE_3868 16'h3802
`define TANH_LUT_POSITIVE_3870 16'h3808
`define TANH_LUT_POSITIVE_3878 16'h380E
`define TANH_LUT_POSITIVE_3880 16'h3814
`define TANH_LUT_POSITIVE_3888 16'h381A
`define TANH_LUT_POSITIVE_3890 16'h3820
`define TANH_LUT_POSITIVE_3898 16'h3826
`define TANH_LUT_POSITIVE_38A0 16'h382C
`define TANH_LUT_POSITIVE_38A8 16'h3831
`define TANH_LUT_POSITIVE_38B0 16'h3837
`define TANH_LUT_POSITIVE_38B8 16'h383D
`define TANH_LUT_POSITIVE_38C0 16'h3843
`define TANH_LUT_POSITIVE_38C8 16'h3848
`define TANH_LUT_POSITIVE_38D0 16'h384E
`define TANH_LUT_POSITIVE_38D8 16'h3854
`define TANH_LUT_POSITIVE_38E0 16'h3859
`define TANH_LUT_POSITIVE_38E8 16'h385F
`define TANH_LUT_POSITIVE_38F0 16'h3865
`define TANH_LUT_POSITIVE_38F8 16'h386A
`define TANH_LUT_POSITIVE_3900 16'h3870
`define TANH_LUT_POSITIVE_3908 16'h3875
`define TANH_LUT_POSITIVE_3910 16'h387B
`define TANH_LUT_POSITIVE_3918 16'h3880
`define TANH_LUT_POSITIVE_3920 16'h3886
`define TANH_LUT_POSITIVE_3928 16'h388B
`define TANH_LUT_POSITIVE_3930 16'h3891
`define TANH_LUT_POSITIVE_3938 16'h3896
`define TANH_LUT_POSITIVE_3940 16'h389B
`define TANH_LUT_POSITIVE_3948 16'h38A1
`define TANH_LUT_POSITIVE_3950 16'h38A6
`define TANH_LUT_POSITIVE_3958 16'h38AB
`define TANH_LUT_POSITIVE_3960 16'h38B1
`define TANH_LUT_POSITIVE_3968 16'h38B6
`define TANH_LUT_POSITIVE_3970 16'h38BB
`define TANH_LUT_POSITIVE_3978 16'h38C0
`define TANH_LUT_POSITIVE_3980 16'h38C5
`define TANH_LUT_POSITIVE_3988 16'h38CB
`define TANH_LUT_POSITIVE_3990 16'h38D0
`define TANH_LUT_POSITIVE_3998 16'h38D5
`define TANH_LUT_POSITIVE_39A0 16'h38DA
`define TANH_LUT_POSITIVE_39A8 16'h38DF
`define TANH_LUT_POSITIVE_39B0 16'h38E4
`define TANH_LUT_POSITIVE_39B8 16'h38E9
`define TANH_LUT_POSITIVE_39C0 16'h38EE
`define TANH_LUT_POSITIVE_39C8 16'h38F3
`define TANH_LUT_POSITIVE_39D0 16'h38F8
`define TANH_LUT_POSITIVE_39D8 16'h38FD
`define TANH_LUT_POSITIVE_39E0 16'h3902
`define TANH_LUT_POSITIVE_39E8 16'h3906
`define TANH_LUT_POSITIVE_39F0 16'h390B
`define TANH_LUT_POSITIVE_39F8 16'h3910
`define TANH_LUT_POSITIVE_3A00 16'h3915
`define TANH_LUT_POSITIVE_3A08 16'h391A
`define TANH_LUT_POSITIVE_3A10 16'h391E
`define TANH_LUT_POSITIVE_3A18 16'h3923
`define TANH_LUT_POSITIVE_3A20 16'h3928
`define TANH_LUT_POSITIVE_3A28 16'h392C
`define TANH_LUT_POSITIVE_3A30 16'h3931
`define TANH_LUT_POSITIVE_3A38 16'h3936
`define TANH_LUT_POSITIVE_3A40 16'h393A
`define TANH_LUT_POSITIVE_3A48 16'h393F
`define TANH_LUT_POSITIVE_3A50 16'h3943
`define TANH_LUT_POSITIVE_3A58 16'h3948
`define TANH_LUT_POSITIVE_3A60 16'h394C
`define TANH_LUT_POSITIVE_3A68 16'h3951
`define TANH_LUT_POSITIVE_3A70 16'h3955
`define TANH_LUT_POSITIVE_3A78 16'h395A
`define TANH_LUT_POSITIVE_3A80 16'h395E
`define TANH_LUT_POSITIVE_3A88 16'h3963
`define TANH_LUT_POSITIVE_3A90 16'h3967
`define TANH_LUT_POSITIVE_3A98 16'h396B
`define TANH_LUT_POSITIVE_3AA0 16'h3970
`define TANH_LUT_POSITIVE_3AA8 16'h3974
`define TANH_LUT_POSITIVE_3AB0 16'h3978
`define TANH_LUT_POSITIVE_3AB8 16'h397C
`define TANH_LUT_POSITIVE_3AC0 16'h3981
`define TANH_LUT_POSITIVE_3AC8 16'h3985
`define TANH_LUT_POSITIVE_3AD0 16'h3989
`define TANH_LUT_POSITIVE_3AD8 16'h398D
`define TANH_LUT_POSITIVE_3AE0 16'h3991
`define TANH_LUT_POSITIVE_3AE8 16'h3995
`define TANH_LUT_POSITIVE_3AF0 16'h3999
`define TANH_LUT_POSITIVE_3AF8 16'h399E
`define TANH_LUT_POSITIVE_3B00 16'h39A2
`define TANH_LUT_POSITIVE_3B08 16'h39A6
`define TANH_LUT_POSITIVE_3B10 16'h39AA
`define TANH_LUT_POSITIVE_3B18 16'h39AE
`define TANH_LUT_POSITIVE_3B20 16'h39B2
`define TANH_LUT_POSITIVE_3B28 16'h39B6
`define TANH_LUT_POSITIVE_3B30 16'h39B9
`define TANH_LUT_POSITIVE_3B38 16'h39BD
`define TANH_LUT_POSITIVE_3B40 16'h39C1
`define TANH_LUT_POSITIVE_3B48 16'h39C5
`define TANH_LUT_POSITIVE_3B50 16'h39C9
`define TANH_LUT_POSITIVE_3B58 16'h39CD
`define TANH_LUT_POSITIVE_3B60 16'h39D0
`define TANH_LUT_POSITIVE_3B68 16'h39D4
`define TANH_LUT_POSITIVE_3B70 16'h39D8
`define TANH_LUT_POSITIVE_3B78 16'h39DC
`define TANH_LUT_POSITIVE_3B80 16'h39DF
`define TANH_LUT_POSITIVE_3B88 16'h39E3
`define TANH_LUT_POSITIVE_3B90 16'h39E7
`define TANH_LUT_POSITIVE_3B98 16'h39EA
`define TANH_LUT_POSITIVE_3BA0 16'h39EE
`define TANH_LUT_POSITIVE_3BA8 16'h39F2
`define TANH_LUT_POSITIVE_3BB0 16'h39F5
`define TANH_LUT_POSITIVE_3BB8 16'h39F9
`define TANH_LUT_POSITIVE_3BC0 16'h39FC
`define TANH_LUT_POSITIVE_3BC8 16'h3A00
`define TANH_LUT_POSITIVE_3BD0 16'h3A03
`define TANH_LUT_POSITIVE_3BD8 16'h3A07
`define TANH_LUT_POSITIVE_3BE0 16'h3A0A
`define TANH_LUT_POSITIVE_3BE8 16'h3A0E
`define TANH_LUT_POSITIVE_3BF0 16'h3A11
`define TANH_LUT_POSITIVE_3BF8 16'h3A14
`define TANH_LUT_POSITIVE_3C00 16'h3A18
`define TANH_LUT_POSITIVE_3C08 16'h3A1E
`define TANH_LUT_POSITIVE_3C10 16'h3A25
`define TANH_LUT_POSITIVE_3C18 16'h3A2C
`define TANH_LUT_POSITIVE_3C20 16'h3A32
`define TANH_LUT_POSITIVE_3C28 16'h3A38
`define TANH_LUT_POSITIVE_3C30 16'h3A3F
`define TANH_LUT_POSITIVE_3C38 16'h3A45
`define TANH_LUT_POSITIVE_3C40 16'h3A4B
`define TANH_LUT_POSITIVE_3C48 16'h3A51
`define TANH_LUT_POSITIVE_3C50 16'h3A57
`define TANH_LUT_POSITIVE_3C58 16'h3A5D
`define TANH_LUT_POSITIVE_3C60 16'h3A63
`define TANH_LUT_POSITIVE_3C68 16'h3A69
`define TANH_LUT_POSITIVE_3C70 16'h3A6E
`define TANH_LUT_POSITIVE_3C78 16'h3A74
`define TANH_LUT_POSITIVE_3C80 16'h3A79
`define TANH_LUT_POSITIVE_3C88 16'h3A7F
`define TANH_LUT_POSITIVE_3C90 16'h3A84
`define TANH_LUT_POSITIVE_3C98 16'h3A8A
`define TANH_LUT_POSITIVE_3CA0 16'h3A8F
`define TANH_LUT_POSITIVE_3CA8 16'h3A94
`define TANH_LUT_POSITIVE_3CB0 16'h3A99
`define TANH_LUT_POSITIVE_3CB8 16'h3A9E
`define TANH_LUT_POSITIVE_3CC0 16'h3AA3
`define TANH_LUT_POSITIVE_3CC8 16'h3AA8
`define TANH_LUT_POSITIVE_3CD0 16'h3AAD
`define TANH_LUT_POSITIVE_3CD8 16'h3AB2
`define TANH_LUT_POSITIVE_3CE0 16'h3AB7
`define TANH_LUT_POSITIVE_3CE8 16'h3ABC
`define TANH_LUT_POSITIVE_3CF0 16'h3AC0
`define TANH_LUT_POSITIVE_3CF8 16'h3AC5
`define TANH_LUT_POSITIVE_3D00 16'h3AC9
`define TANH_LUT_POSITIVE_3D08 16'h3ACE
`define TANH_LUT_POSITIVE_3D10 16'h3AD2
`define TANH_LUT_POSITIVE_3D18 16'h3AD6
`define TANH_LUT_POSITIVE_3D20 16'h3ADB
`define TANH_LUT_POSITIVE_3D28 16'h3ADF
`define TANH_LUT_POSITIVE_3D30 16'h3AE3
`define TANH_LUT_POSITIVE_3D38 16'h3AE7
`define TANH_LUT_POSITIVE_3D40 16'h3AEB
`define TANH_LUT_POSITIVE_3D48 16'h3AEF
`define TANH_LUT_POSITIVE_3D50 16'h3AF3
`define TANH_LUT_POSITIVE_3D58 16'h3AF7
`define TANH_LUT_POSITIVE_3D60 16'h3AFB
`define TANH_LUT_POSITIVE_3D68 16'h3AFF
`define TANH_LUT_POSITIVE_3D70 16'h3B03
`define TANH_LUT_POSITIVE_3D78 16'h3B06
`define TANH_LUT_POSITIVE_3D80 16'h3B0A
`define TANH_LUT_POSITIVE_3D88 16'h3B0D
`define TANH_LUT_POSITIVE_3D90 16'h3B11
`define TANH_LUT_POSITIVE_3D98 16'h3B15
`define TANH_LUT_POSITIVE_3DA0 16'h3B18
`define TANH_LUT_POSITIVE_3DA8 16'h3B1B
`define TANH_LUT_POSITIVE_3DB0 16'h3B1F
`define TANH_LUT_POSITIVE_3DB8 16'h3B22
`define TANH_LUT_POSITIVE_3DC0 16'h3B25
`define TANH_LUT_POSITIVE_3DC8 16'h3B28
`define TANH_LUT_POSITIVE_3DD0 16'h3B2C
`define TANH_LUT_POSITIVE_3DD8 16'h3B2F
`define TANH_LUT_POSITIVE_3DE0 16'h3B32
`define TANH_LUT_POSITIVE_3DE8 16'h3B35
`define TANH_LUT_POSITIVE_3DF0 16'h3B38
`define TANH_LUT_POSITIVE_3DF8 16'h3B3B
`define TANH_LUT_POSITIVE_3E00 16'h3B3E
`define TANH_LUT_POSITIVE_3E08 16'h3B41
`define TANH_LUT_POSITIVE_3E10 16'h3B43
`define TANH_LUT_POSITIVE_3E18 16'h3B46
`define TANH_LUT_POSITIVE_3E20 16'h3B49
`define TANH_LUT_POSITIVE_3E28 16'h3B4C
`define TANH_LUT_POSITIVE_3E30 16'h3B4E
`define TANH_LUT_POSITIVE_3E38 16'h3B51
`define TANH_LUT_POSITIVE_3E40 16'h3B54
`define TANH_LUT_POSITIVE_3E48 16'h3B56
`define TANH_LUT_POSITIVE_3E50 16'h3B59
`define TANH_LUT_POSITIVE_3E58 16'h3B5B
`define TANH_LUT_POSITIVE_3E60 16'h3B5E
`define TANH_LUT_POSITIVE_3E68 16'h3B60
`define TANH_LUT_POSITIVE_3E70 16'h3B62
`define TANH_LUT_POSITIVE_3E78 16'h3B65
`define TANH_LUT_POSITIVE_3E80 16'h3B67
`define TANH_LUT_POSITIVE_3E88 16'h3B69
`define TANH_LUT_POSITIVE_3E90 16'h3B6C
`define TANH_LUT_POSITIVE_3E98 16'h3B6E
`define TANH_LUT_POSITIVE_3EA0 16'h3B70
`define TANH_LUT_POSITIVE_3EA8 16'h3B72
`define TANH_LUT_POSITIVE_3EB0 16'h3B74
`define TANH_LUT_POSITIVE_3EB8 16'h3B76
`define TANH_LUT_POSITIVE_3EC0 16'h3B78
`define TANH_LUT_POSITIVE_3EC8 16'h3B7B
`define TANH_LUT_POSITIVE_3ED0 16'h3B7D
`define TANH_LUT_POSITIVE_3ED8 16'h3B7E
`define TANH_LUT_POSITIVE_3EE0 16'h3B80
`define TANH_LUT_POSITIVE_3EE8 16'h3B82
`define TANH_LUT_POSITIVE_3EF0 16'h3B84
`define TANH_LUT_POSITIVE_3EF8 16'h3B86
`define TANH_LUT_POSITIVE_3F00 16'h3B88
`define TANH_LUT_POSITIVE_3F08 16'h3B8A
`define TANH_LUT_POSITIVE_3F10 16'h3B8C
`define TANH_LUT_POSITIVE_3F18 16'h3B8D
`define TANH_LUT_POSITIVE_3F20 16'h3B8F
`define TANH_LUT_POSITIVE_3F28 16'h3B91
`define TANH_LUT_POSITIVE_3F30 16'h3B92
`define TANH_LUT_POSITIVE_3F38 16'h3B94
`define TANH_LUT_POSITIVE_3F40 16'h3B96
`define TANH_LUT_POSITIVE_3F48 16'h3B97
`define TANH_LUT_POSITIVE_3F50 16'h3B99
`define TANH_LUT_POSITIVE_3F58 16'h3B9A
`define TANH_LUT_POSITIVE_3F60 16'h3B9C
`define TANH_LUT_POSITIVE_3F68 16'h3B9D
`define TANH_LUT_POSITIVE_3F70 16'h3B9F
`define TANH_LUT_POSITIVE_3F78 16'h3BA0
`define TANH_LUT_POSITIVE_3F80 16'h3BA2
`define TANH_LUT_POSITIVE_3F88 16'h3BA3
`define TANH_LUT_POSITIVE_3F90 16'h3BA5
`define TANH_LUT_POSITIVE_3F98 16'h3BA6
`define TANH_LUT_POSITIVE_3FA0 16'h3BA7
`define TANH_LUT_POSITIVE_3FA8 16'h3BA9
`define TANH_LUT_POSITIVE_3FB0 16'h3BAA
`define TANH_LUT_POSITIVE_3FB8 16'h3BAB
`define TANH_LUT_POSITIVE_3FC0 16'h3BAD
`define TANH_LUT_POSITIVE_3FC8 16'h3BAE
`define TANH_LUT_POSITIVE_3FD0 16'h3BAF
`define TANH_LUT_POSITIVE_3FD8 16'h3BB0
`define TANH_LUT_POSITIVE_3FE0 16'h3BB2
`define TANH_LUT_POSITIVE_3FE8 16'h3BB3
`define TANH_LUT_POSITIVE_3FF0 16'h3BB4
`define TANH_LUT_POSITIVE_3FF8 16'h3BB5
`define TANH_LUT_POSITIVE_4000 16'h3BB6
`define TANH_LUT_POSITIVE_4008 16'h3BB9
`define TANH_LUT_POSITIVE_4010 16'h3BBB
`define TANH_LUT_POSITIVE_4018 16'h3BBD
`define TANH_LUT_POSITIVE_4020 16'h3BBF
`define TANH_LUT_POSITIVE_4028 16'h3BC1
`define TANH_LUT_POSITIVE_4030 16'h3BC3
`define TANH_LUT_POSITIVE_4038 16'h3BC5
`define TANH_LUT_POSITIVE_4040 16'h3BC6
`define TANH_LUT_POSITIVE_4048 16'h3BC8
`define TANH_LUT_POSITIVE_4050 16'h3BCA
`define TANH_LUT_POSITIVE_4058 16'h3BCB
`define TANH_LUT_POSITIVE_4060 16'h3BCD
`define TANH_LUT_POSITIVE_4068 16'h3BCF
`define TANH_LUT_POSITIVE_4070 16'h3BD0
`define TANH_LUT_POSITIVE_4078 16'h3BD2
`define TANH_LUT_POSITIVE_4080 16'h3BD3
`define TANH_LUT_POSITIVE_4088 16'h3BD4
`define TANH_LUT_POSITIVE_4090 16'h3BD6
`define TANH_LUT_POSITIVE_4098 16'h3BD7
`define TANH_LUT_POSITIVE_40A0 16'h3BD8
`define TANH_LUT_POSITIVE_40A8 16'h3BD9
`define TANH_LUT_POSITIVE_40B0 16'h3BDB
`define TANH_LUT_POSITIVE_40B8 16'h3BDC
`define TANH_LUT_POSITIVE_40C0 16'h3BDD
`define TANH_LUT_POSITIVE_40C8 16'h3BDE
`define TANH_LUT_POSITIVE_40D0 16'h3BDF
`define TANH_LUT_POSITIVE_40D8 16'h3BE0
`define TANH_LUT_POSITIVE_40E0 16'h3BE1
`define TANH_LUT_POSITIVE_40E8 16'h3BE2
`define TANH_LUT_POSITIVE_40F0 16'h3BE3
`define TANH_LUT_POSITIVE_40F8 16'h3BE4
`define TANH_LUT_POSITIVE_4100 16'h3BE5
`define TANH_LUT_POSITIVE_4108 16'h3BE5
`define TANH_LUT_POSITIVE_4110 16'h3BE6
`define TANH_LUT_POSITIVE_4118 16'h3BE7
`define TANH_LUT_POSITIVE_4120 16'h3BE8
`define TANH_LUT_POSITIVE_4128 16'h3BE9
`define TANH_LUT_POSITIVE_4130 16'h3BE9
`define TANH_LUT_POSITIVE_4138 16'h3BEA
`define TANH_LUT_POSITIVE_4140 16'h3BEB
`define TANH_LUT_POSITIVE_4148 16'h3BEB
`define TANH_LUT_POSITIVE_4150 16'h3BEC
`define TANH_LUT_POSITIVE_4158 16'h3BED
`define TANH_LUT_POSITIVE_4160 16'h3BED
`define TANH_LUT_POSITIVE_4168 16'h3BEE
`define TANH_LUT_POSITIVE_4170 16'h3BEE
`define TANH_LUT_POSITIVE_4178 16'h3BEF
`define TANH_LUT_POSITIVE_4180 16'h3BEF
`define TANH_LUT_POSITIVE_4188 16'h3BF0
`define TANH_LUT_POSITIVE_4190 16'h3BF0
`define TANH_LUT_POSITIVE_4198 16'h3BF1
`define TANH_LUT_POSITIVE_41A0 16'h3BF1
`define TANH_LUT_POSITIVE_41A8 16'h3BF2
`define TANH_LUT_POSITIVE_41B0 16'h3BF2
`define TANH_LUT_POSITIVE_41B8 16'h3BF3
`define TANH_LUT_POSITIVE_41C0 16'h3BF3
`define TANH_LUT_POSITIVE_41C8 16'h3BF3
`define TANH_LUT_POSITIVE_41D0 16'h3BF4
`define TANH_LUT_POSITIVE_41D8 16'h3BF4
`define TANH_LUT_POSITIVE_41E0 16'h3BF5
`define TANH_LUT_POSITIVE_41E8 16'h3BF5
`define TANH_LUT_POSITIVE_41F0 16'h3BF5
`define TANH_LUT_POSITIVE_41F8 16'h3BF6
`define TANH_LUT_POSITIVE_4200 16'h3BF6
`define TANH_LUT_POSITIVE_4208 16'h3BF6
`define TANH_LUT_POSITIVE_4210 16'h3BF6
`define TANH_LUT_POSITIVE_4218 16'h3BF7
`define TANH_LUT_POSITIVE_4220 16'h3BF7
`define TANH_LUT_POSITIVE_4228 16'h3BF7
`define TANH_LUT_POSITIVE_4230 16'h3BF8
`define TANH_LUT_POSITIVE_4238 16'h3BF8
`define TANH_LUT_POSITIVE_4240 16'h3BF8
`define TANH_LUT_POSITIVE_4248 16'h3BF8
`define TANH_LUT_POSITIVE_4250 16'h3BF9
`define TANH_LUT_POSITIVE_4258 16'h3BF9
`define TANH_LUT_POSITIVE_4260 16'h3BF9
`define TANH_LUT_POSITIVE_4268 16'h3BF9
`define TANH_LUT_POSITIVE_4270 16'h3BF9
`define TANH_LUT_POSITIVE_4278 16'h3BFA
`define TANH_LUT_POSITIVE_4280 16'h3BFA
`define TANH_LUT_POSITIVE_4288 16'h3BFA
`define TANH_LUT_POSITIVE_4290 16'h3BFA
`define TANH_LUT_POSITIVE_4298 16'h3BFA
`define TANH_LUT_POSITIVE_42A0 16'h3BFB
`define TANH_LUT_POSITIVE_42A8 16'h3BFB
`define TANH_LUT_POSITIVE_42B0 16'h3BFB
`define TANH_LUT_POSITIVE_42B8 16'h3BFB
`define TANH_LUT_POSITIVE_42C0 16'h3BFB
`define TANH_LUT_POSITIVE_42C8 16'h3BFB
`define TANH_LUT_POSITIVE_42D0 16'h3BFB
`define TANH_LUT_POSITIVE_42D8 16'h3BFC
