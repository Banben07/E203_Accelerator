`define CUBE_LUT_2745 16'h2744
`define CUBE_LUT_2746 16'h2745
`define CUBE_LUT_2747 16'h2746
`define CUBE_LUT_2748 16'h2747
`define CUBE_LUT_2749 16'h2748
`define CUBE_LUT_274A 16'h2749
`define CUBE_LUT_274B 16'h274A
`define CUBE_LUT_274C 16'h274B
`define CUBE_LUT_274D 16'h274C
`define CUBE_LUT_274E 16'h274D
`define CUBE_LUT_274F 16'h274E
`define CUBE_LUT_2750 16'h274F
`define CUBE_LUT_2751 16'h2750
`define CUBE_LUT_2752 16'h2751
`define CUBE_LUT_2753 16'h2752
`define CUBE_LUT_2754 16'h2753
`define CUBE_LUT_2755 16'h2754
`define CUBE_LUT_2756 16'h2755
`define CUBE_LUT_2757 16'h2756
`define CUBE_LUT_2758 16'h2757
`define CUBE_LUT_2759 16'h2758
`define CUBE_LUT_275A 16'h2759
`define CUBE_LUT_275B 16'h275A
`define CUBE_LUT_275C 16'h275B
`define CUBE_LUT_275D 16'h275C
`define CUBE_LUT_275E 16'h275D
`define CUBE_LUT_275F 16'h275E
`define CUBE_LUT_2760 16'h275F
`define CUBE_LUT_2761 16'h2760
`define CUBE_LUT_2762 16'h2761
`define CUBE_LUT_2763 16'h2762
`define CUBE_LUT_2764 16'h2763
`define CUBE_LUT_2765 16'h2764
`define CUBE_LUT_2766 16'h2765
`define CUBE_LUT_2767 16'h2766
`define CUBE_LUT_2768 16'h2767
`define CUBE_LUT_2769 16'h2768
`define CUBE_LUT_276A 16'h2769
`define CUBE_LUT_276B 16'h276A
`define CUBE_LUT_276C 16'h276B
`define CUBE_LUT_276D 16'h276C
`define CUBE_LUT_276E 16'h276D
`define CUBE_LUT_276F 16'h276E
`define CUBE_LUT_2770 16'h276F
`define CUBE_LUT_2771 16'h2770
`define CUBE_LUT_2772 16'h2771
`define CUBE_LUT_2773 16'h2772
`define CUBE_LUT_2774 16'h2773
`define CUBE_LUT_2775 16'h2774
`define CUBE_LUT_2776 16'h2775
`define CUBE_LUT_2777 16'h2776
`define CUBE_LUT_2778 16'h2777
`define CUBE_LUT_2779 16'h2778
`define CUBE_LUT_277A 16'h2779
`define CUBE_LUT_277B 16'h277A
`define CUBE_LUT_277C 16'h277B
`define CUBE_LUT_277D 16'h277C
`define CUBE_LUT_277E 16'h277D
`define CUBE_LUT_277F 16'h277E
`define CUBE_LUT_2780 16'h277F
`define CUBE_LUT_2781 16'h2780
`define CUBE_LUT_2782 16'h2781
`define CUBE_LUT_2783 16'h2782
`define CUBE_LUT_2784 16'h2783
`define CUBE_LUT_2785 16'h2784
`define CUBE_LUT_2786 16'h2785
`define CUBE_LUT_2787 16'h2786
`define CUBE_LUT_2788 16'h2787
`define CUBE_LUT_2789 16'h2788
`define CUBE_LUT_278A 16'h2789
`define CUBE_LUT_278B 16'h278A
`define CUBE_LUT_278C 16'h278B
`define CUBE_LUT_278D 16'h278C
`define CUBE_LUT_278E 16'h278D
`define CUBE_LUT_278F 16'h278E
`define CUBE_LUT_2790 16'h278F
`define CUBE_LUT_2791 16'h2790
`define CUBE_LUT_2792 16'h2791
`define CUBE_LUT_2793 16'h2792
`define CUBE_LUT_2794 16'h2793
`define CUBE_LUT_2795 16'h2794
`define CUBE_LUT_2796 16'h2795
`define CUBE_LUT_2797 16'h2796
`define CUBE_LUT_2798 16'h2797
`define CUBE_LUT_2799 16'h2798
`define CUBE_LUT_279A 16'h2799
`define CUBE_LUT_279B 16'h279A
`define CUBE_LUT_279C 16'h279B
`define CUBE_LUT_279D 16'h279C
`define CUBE_LUT_279E 16'h279D
`define CUBE_LUT_279F 16'h279E
`define CUBE_LUT_27A0 16'h279F
`define CUBE_LUT_27A1 16'h27A0
`define CUBE_LUT_27A2 16'h27A1
`define CUBE_LUT_27A3 16'h27A2
`define CUBE_LUT_27A4 16'h27A3
`define CUBE_LUT_27A5 16'h27A4
`define CUBE_LUT_27A6 16'h27A5
`define CUBE_LUT_27A7 16'h27A6
`define CUBE_LUT_27A8 16'h27A7
`define CUBE_LUT_27A9 16'h27A8
`define CUBE_LUT_27AA 16'h27A9
`define CUBE_LUT_27AB 16'h27AA
`define CUBE_LUT_27AC 16'h27AB
`define CUBE_LUT_27AD 16'h27AC
`define CUBE_LUT_27AE 16'h27AD
`define CUBE_LUT_27AF 16'h27AE
`define CUBE_LUT_27B0 16'h27AF
`define CUBE_LUT_27B1 16'h27B0
`define CUBE_LUT_27B2 16'h27B1
`define CUBE_LUT_27B3 16'h27B2
`define CUBE_LUT_27B4 16'h27B3
`define CUBE_LUT_27B5 16'h27B4
`define CUBE_LUT_27B6 16'h27B5
`define CUBE_LUT_27B7 16'h27B6
`define CUBE_LUT_27B8 16'h27B7
`define CUBE_LUT_27B9 16'h27B8
`define CUBE_LUT_27BA 16'h27B9
`define CUBE_LUT_27BB 16'h27BA
`define CUBE_LUT_27BC 16'h27BB
`define CUBE_LUT_27BD 16'h27BC
`define CUBE_LUT_27BE 16'h27BD
`define CUBE_LUT_27BF 16'h27BE
`define CUBE_LUT_27C0 16'h27BF
`define CUBE_LUT_27C1 16'h27C0
`define CUBE_LUT_27C2 16'h27C1
`define CUBE_LUT_27C3 16'h27C2
`define CUBE_LUT_27C4 16'h27C3
`define CUBE_LUT_27C5 16'h27C4
`define CUBE_LUT_27C6 16'h27C5
`define CUBE_LUT_27C7 16'h27C6
`define CUBE_LUT_27C8 16'h27C7
`define CUBE_LUT_27C9 16'h27C8
`define CUBE_LUT_27CA 16'h27C9
`define CUBE_LUT_27CB 16'h27CA
`define CUBE_LUT_27CC 16'h27CB
`define CUBE_LUT_27CD 16'h27CC
`define CUBE_LUT_27CE 16'h27CD
`define CUBE_LUT_27CF 16'h27CE
`define CUBE_LUT_27D0 16'h27CF
`define CUBE_LUT_27D1 16'h27D0
`define CUBE_LUT_27D2 16'h27D1
`define CUBE_LUT_27D3 16'h27D2
`define CUBE_LUT_27D4 16'h27D3
`define CUBE_LUT_27D5 16'h27D4
`define CUBE_LUT_27D6 16'h27D5
`define CUBE_LUT_27D7 16'h27D6
`define CUBE_LUT_27D8 16'h27D7
`define CUBE_LUT_27D9 16'h27D8
`define CUBE_LUT_27DA 16'h27D9
`define CUBE_LUT_27DB 16'h27DA
`define CUBE_LUT_27DC 16'h27DB
`define CUBE_LUT_27DD 16'h27DC
`define CUBE_LUT_27DE 16'h27DD
`define CUBE_LUT_27DF 16'h27DE
`define CUBE_LUT_27E0 16'h27DF
`define CUBE_LUT_27E1 16'h27E0
`define CUBE_LUT_27E2 16'h27E1
`define CUBE_LUT_27E3 16'h27E2
`define CUBE_LUT_27E4 16'h27E3
`define CUBE_LUT_27E5 16'h27E4
`define CUBE_LUT_27E6 16'h27E5
`define CUBE_LUT_27E7 16'h27E6
`define CUBE_LUT_27E8 16'h27E7
`define CUBE_LUT_27E9 16'h27E8
`define CUBE_LUT_27EA 16'h27E9
`define CUBE_LUT_27EB 16'h27EA
`define CUBE_LUT_27EC 16'h27EB
`define CUBE_LUT_27ED 16'h27EC
`define CUBE_LUT_27EE 16'h27ED
`define CUBE_LUT_27EF 16'h27EE
`define CUBE_LUT_27F0 16'h27EF
`define CUBE_LUT_27F1 16'h27F0
`define CUBE_LUT_27F2 16'h27F1
`define CUBE_LUT_27F3 16'h27F2
`define CUBE_LUT_27F4 16'h27F3
`define CUBE_LUT_27F5 16'h27F4
`define CUBE_LUT_27F6 16'h27F5
`define CUBE_LUT_27F7 16'h27F6
`define CUBE_LUT_27F8 16'h27F7
`define CUBE_LUT_27F9 16'h27F8
`define CUBE_LUT_27FA 16'h27F9
`define CUBE_LUT_27FB 16'h27FA
`define CUBE_LUT_27FC 16'h27FB
`define CUBE_LUT_27FD 16'h27FC
`define CUBE_LUT_27FE 16'h27FD
`define CUBE_LUT_27FF 16'h27FE
`define CUBE_LUT_2800 16'h27FF

`define CUBE_LUT_2801 16'h2801
`define CUBE_LUT_2802 16'h2802
`define CUBE_LUT_2803 16'h2803
`define CUBE_LUT_2804 16'h2804
`define CUBE_LUT_2805 16'h2805
`define CUBE_LUT_2806 16'h2806
`define CUBE_LUT_2807 16'h2807
`define CUBE_LUT_2808 16'h2808
`define CUBE_LUT_2809 16'h2809
`define CUBE_LUT_280A 16'h280A
`define CUBE_LUT_280B 16'h280B
`define CUBE_LUT_280C 16'h280C
`define CUBE_LUT_280D 16'h280D
`define CUBE_LUT_280E 16'h280E
`define CUBE_LUT_280F 16'h280F
`define CUBE_LUT_2810 16'h2810
`define CUBE_LUT_2811 16'h2811
`define CUBE_LUT_2812 16'h2812
`define CUBE_LUT_2813 16'h2813
`define CUBE_LUT_2814 16'h2814
`define CUBE_LUT_2815 16'h2815
`define CUBE_LUT_2816 16'h2816
`define CUBE_LUT_2817 16'h2817
`define CUBE_LUT_2818 16'h2818
`define CUBE_LUT_2819 16'h2819
`define CUBE_LUT_281A 16'h281A
`define CUBE_LUT_281B 16'h281B
`define CUBE_LUT_281C 16'h281C
`define CUBE_LUT_281D 16'h281D
`define CUBE_LUT_281E 16'h281E
`define CUBE_LUT_281F 16'h281F
`define CUBE_LUT_2820 16'h2820
`define CUBE_LUT_2821 16'h2821
`define CUBE_LUT_2822 16'h2822
`define CUBE_LUT_2823 16'h2823
`define CUBE_LUT_2824 16'h2824
`define CUBE_LUT_2825 16'h2825
`define CUBE_LUT_2826 16'h2826
`define CUBE_LUT_2827 16'h2827
`define CUBE_LUT_2828 16'h2828
`define CUBE_LUT_2829 16'h2829
`define CUBE_LUT_282A 16'h282A
`define CUBE_LUT_282B 16'h282B
`define CUBE_LUT_282C 16'h282C
`define CUBE_LUT_282D 16'h282D
`define CUBE_LUT_282E 16'h282E
`define CUBE_LUT_282F 16'h282F
`define CUBE_LUT_2830 16'h2830
`define CUBE_LUT_2831 16'h2831
`define CUBE_LUT_2832 16'h2832
`define CUBE_LUT_2833 16'h2833
`define CUBE_LUT_2834 16'h2834
`define CUBE_LUT_2835 16'h2835
`define CUBE_LUT_2836 16'h2836
`define CUBE_LUT_2837 16'h2837
`define CUBE_LUT_2838 16'h2838
`define CUBE_LUT_2839 16'h2839
`define CUBE_LUT_283A 16'h283A
`define CUBE_LUT_283B 16'h283B
`define CUBE_LUT_283C 16'h283C
`define CUBE_LUT_283D 16'h283D
`define CUBE_LUT_283E 16'h283E
`define CUBE_LUT_283F 16'h283F
`define CUBE_LUT_2840 16'h2840
`define CUBE_LUT_2841 16'h2841
`define CUBE_LUT_2842 16'h2842
`define CUBE_LUT_2843 16'h2843
`define CUBE_LUT_2844 16'h2844
`define CUBE_LUT_2845 16'h2845
`define CUBE_LUT_2846 16'h2846
`define CUBE_LUT_2847 16'h2847
`define CUBE_LUT_2848 16'h2848
`define CUBE_LUT_2849 16'h2849
`define CUBE_LUT_284A 16'h284A
`define CUBE_LUT_284B 16'h284B
`define CUBE_LUT_284C 16'h284C
`define CUBE_LUT_284D 16'h284D
`define CUBE_LUT_284E 16'h284E
`define CUBE_LUT_284F 16'h284F
`define CUBE_LUT_2850 16'h2850
`define CUBE_LUT_2851 16'h2851
`define CUBE_LUT_2852 16'h2852
`define CUBE_LUT_2853 16'h2853
`define CUBE_LUT_2854 16'h2854
`define CUBE_LUT_2855 16'h2855
`define CUBE_LUT_2856 16'h2856
`define CUBE_LUT_2857 16'h2857
`define CUBE_LUT_2858 16'h2858
`define CUBE_LUT_2859 16'h2859
`define CUBE_LUT_285A 16'h285A
`define CUBE_LUT_285B 16'h285B
`define CUBE_LUT_285C 16'h285C
`define CUBE_LUT_285D 16'h285D
`define CUBE_LUT_285E 16'h285E
`define CUBE_LUT_285F 16'h285F
`define CUBE_LUT_2860 16'h2860
`define CUBE_LUT_2861 16'h2861
`define CUBE_LUT_2862 16'h2862
`define CUBE_LUT_2863 16'h2863
`define CUBE_LUT_2864 16'h2864
`define CUBE_LUT_2865 16'h2865
`define CUBE_LUT_2866 16'h2866
`define CUBE_LUT_2867 16'h2867
`define CUBE_LUT_2868 16'h2868
`define CUBE_LUT_2869 16'h2869
`define CUBE_LUT_286A 16'h286A
`define CUBE_LUT_286B 16'h286B
`define CUBE_LUT_286C 16'h286C
`define CUBE_LUT_286D 16'h286D
`define CUBE_LUT_286E 16'h286E
`define CUBE_LUT_286F 16'h286F
`define CUBE_LUT_2870 16'h2870
`define CUBE_LUT_2871 16'h2871
`define CUBE_LUT_2872 16'h2872
`define CUBE_LUT_2873 16'h2873
`define CUBE_LUT_2874 16'h2874
`define CUBE_LUT_2875 16'h2875
`define CUBE_LUT_2876 16'h2876
`define CUBE_LUT_2877 16'h2877
`define CUBE_LUT_2878 16'h2878
`define CUBE_LUT_2879 16'h2879
`define CUBE_LUT_287A 16'h287A
`define CUBE_LUT_287B 16'h287B
`define CUBE_LUT_287C 16'h287C
`define CUBE_LUT_287D 16'h287D
`define CUBE_LUT_287E 16'h287E
`define CUBE_LUT_287F 16'h287F
`define CUBE_LUT_2880 16'h2880
`define CUBE_LUT_2881 16'h2881
`define CUBE_LUT_2882 16'h2882
`define CUBE_LUT_2883 16'h2883
`define CUBE_LUT_2884 16'h2884
`define CUBE_LUT_2885 16'h2885
`define CUBE_LUT_2886 16'h2886
`define CUBE_LUT_2887 16'h2887
`define CUBE_LUT_2888 16'h2888
`define CUBE_LUT_2889 16'h2889
`define CUBE_LUT_288A 16'h288A
`define CUBE_LUT_288B 16'h288B
`define CUBE_LUT_288C 16'h288C
`define CUBE_LUT_288D 16'h288D
`define CUBE_LUT_288E 16'h288E
`define CUBE_LUT_288F 16'h288F
`define CUBE_LUT_2890 16'h2890
`define CUBE_LUT_2891 16'h2891
`define CUBE_LUT_2892 16'h2892
`define CUBE_LUT_2893 16'h2893
`define CUBE_LUT_2894 16'h2894

`define CUBE_LUT_2895 16'h2894
`define CUBE_LUT_2896 16'h2895
`define CUBE_LUT_2897 16'h2896
`define CUBE_LUT_2898 16'h2897
`define CUBE_LUT_2899 16'h2898
`define CUBE_LUT_289A 16'h2899
`define CUBE_LUT_289B 16'h289A
`define CUBE_LUT_289C 16'h289B
`define CUBE_LUT_289D 16'h289C
`define CUBE_LUT_289E 16'h289D
`define CUBE_LUT_289F 16'h289E
`define CUBE_LUT_28A0 16'h289F
`define CUBE_LUT_28A1 16'h28A0
`define CUBE_LUT_28A2 16'h28A1
`define CUBE_LUT_28A3 16'h28A2
`define CUBE_LUT_28A4 16'h28A3
`define CUBE_LUT_28A5 16'h28A4
`define CUBE_LUT_28A6 16'h28A5
`define CUBE_LUT_28A7 16'h28A6
`define CUBE_LUT_28A8 16'h28A7
`define CUBE_LUT_28A9 16'h28A8
`define CUBE_LUT_28AA 16'h28A9
`define CUBE_LUT_28AB 16'h28AA
`define CUBE_LUT_28AC 16'h28AB
`define CUBE_LUT_28AD 16'h28AC
`define CUBE_LUT_28AE 16'h28AD
`define CUBE_LUT_28AF 16'h28AE
`define CUBE_LUT_28B0 16'h28AF
`define CUBE_LUT_28B1 16'h28B0
`define CUBE_LUT_28B2 16'h28B1
`define CUBE_LUT_28B3 16'h28B2
`define CUBE_LUT_28B4 16'h28B3
`define CUBE_LUT_28B5 16'h28B4
`define CUBE_LUT_28B6 16'h28B5
`define CUBE_LUT_28B7 16'h28B6
`define CUBE_LUT_28B8 16'h28B7
`define CUBE_LUT_28B9 16'h28B8
`define CUBE_LUT_28BA 16'h28B9
`define CUBE_LUT_28BB 16'h28BA
`define CUBE_LUT_28BC 16'h28BB
`define CUBE_LUT_28BD 16'h28BC
`define CUBE_LUT_28BE 16'h28BD
`define CUBE_LUT_28BF 16'h28BE
`define CUBE_LUT_28C0 16'h28BF
`define CUBE_LUT_28C1 16'h28C0
`define CUBE_LUT_28C2 16'h28C1
`define CUBE_LUT_28C3 16'h28C2
`define CUBE_LUT_28C4 16'h28C3
`define CUBE_LUT_28C5 16'h28C4
`define CUBE_LUT_28C6 16'h28C5
`define CUBE_LUT_28C7 16'h28C6
`define CUBE_LUT_28C8 16'h28C7
`define CUBE_LUT_28C9 16'h28C8
`define CUBE_LUT_28CA 16'h28C9
`define CUBE_LUT_28CB 16'h28CA
`define CUBE_LUT_28CC 16'h28CB
`define CUBE_LUT_28CD 16'h28CC
`define CUBE_LUT_28CE 16'h28CD
`define CUBE_LUT_28CF 16'h28CE
`define CUBE_LUT_28D0 16'h28CF
`define CUBE_LUT_28D1 16'h28D0
`define CUBE_LUT_28D2 16'h28D1
`define CUBE_LUT_28D3 16'h28D2
`define CUBE_LUT_28D4 16'h28D3
`define CUBE_LUT_28D5 16'h28D4
`define CUBE_LUT_28D6 16'h28D5
`define CUBE_LUT_28D7 16'h28D6
`define CUBE_LUT_28D8 16'h28D7
`define CUBE_LUT_28D9 16'h28D8
`define CUBE_LUT_28DA 16'h28D9
`define CUBE_LUT_28DB 16'h28DA
`define CUBE_LUT_28DC 16'h28DB
`define CUBE_LUT_28DD 16'h28DC
`define CUBE_LUT_28DE 16'h28DD
`define CUBE_LUT_28DF 16'h28DE
`define CUBE_LUT_28E0 16'h28DF
`define CUBE_LUT_28E1 16'h28E0
`define CUBE_LUT_28E2 16'h28E1
`define CUBE_LUT_28E3 16'h28E2
`define CUBE_LUT_28E4 16'h28E3
`define CUBE_LUT_28E5 16'h28E4
`define CUBE_LUT_28E6 16'h28E5
`define CUBE_LUT_28E7 16'h28E6
`define CUBE_LUT_28E8 16'h28E7
`define CUBE_LUT_28E9 16'h28E8
`define CUBE_LUT_28EA 16'h28E9
`define CUBE_LUT_28EB 16'h28EA
`define CUBE_LUT_28EC 16'h28EB
`define CUBE_LUT_28ED 16'h28EC
`define CUBE_LUT_28EE 16'h28ED
`define CUBE_LUT_28EF 16'h28EE
`define CUBE_LUT_28F0 16'h28EF
`define CUBE_LUT_28F1 16'h28F0
`define CUBE_LUT_28F2 16'h28F1
`define CUBE_LUT_28F3 16'h28F2
`define CUBE_LUT_28F4 16'h28F3
`define CUBE_LUT_28F5 16'h28F4
`define CUBE_LUT_28F6 16'h28F5
`define CUBE_LUT_28F7 16'h28F6
`define CUBE_LUT_28F8 16'h28F7
`define CUBE_LUT_28F9 16'h28F8
`define CUBE_LUT_28FA 16'h28F9
`define CUBE_LUT_28FB 16'h28FA
`define CUBE_LUT_28FC 16'h28FB
`define CUBE_LUT_28FD 16'h28FC
`define CUBE_LUT_28FE 16'h28FD
`define CUBE_LUT_28FF 16'h28FE
`define CUBE_LUT_2900 16'h28FF
`define CUBE_LUT_2901 16'h2900
`define CUBE_LUT_2902 16'h2901
`define CUBE_LUT_2903 16'h2902
`define CUBE_LUT_2904 16'h2903
`define CUBE_LUT_2905 16'h2904
`define CUBE_LUT_2906 16'h2905
`define CUBE_LUT_2907 16'h2906
`define CUBE_LUT_2908 16'h2907
`define CUBE_LUT_2909 16'h2908
`define CUBE_LUT_290A 16'h2909
`define CUBE_LUT_290B 16'h290A
`define CUBE_LUT_290C 16'h290B
`define CUBE_LUT_290D 16'h290C
`define CUBE_LUT_290E 16'h290D
`define CUBE_LUT_290F 16'h290E
`define CUBE_LUT_2910 16'h290F
`define CUBE_LUT_2911 16'h2910
`define CUBE_LUT_2912 16'h2911
`define CUBE_LUT_2913 16'h2912
`define CUBE_LUT_2914 16'h2913
`define CUBE_LUT_2915 16'h2914
`define CUBE_LUT_2916 16'h2915
`define CUBE_LUT_2917 16'h2916
`define CUBE_LUT_2918 16'h2917
`define CUBE_LUT_2919 16'h2918
`define CUBE_LUT_291A 16'h2919
`define CUBE_LUT_291B 16'h291A
`define CUBE_LUT_291C 16'h291B
`define CUBE_LUT_291D 16'h291C
`define CUBE_LUT_291E 16'h291D
`define CUBE_LUT_291F 16'h291E
`define CUBE_LUT_2920 16'h291F
`define CUBE_LUT_2921 16'h2920
`define CUBE_LUT_2922 16'h2921
`define CUBE_LUT_2923 16'h2922
`define CUBE_LUT_2924 16'h2923
`define CUBE_LUT_2925 16'h2924
`define CUBE_LUT_2926 16'h2925
`define CUBE_LUT_2927 16'h2926
`define CUBE_LUT_2928 16'h2927
`define CUBE_LUT_2929 16'h2928
`define CUBE_LUT_292A 16'h2929
`define CUBE_LUT_292B 16'h292A
`define CUBE_LUT_292C 16'h292B
`define CUBE_LUT_292D 16'h292C
`define CUBE_LUT_292E 16'h292D
`define CUBE_LUT_292F 16'h292E
`define CUBE_LUT_2930 16'h292F
`define CUBE_LUT_2931 16'h2930
`define CUBE_LUT_2932 16'h2931
`define CUBE_LUT_2933 16'h2932
`define CUBE_LUT_2934 16'h2933
`define CUBE_LUT_2935 16'h2934
`define CUBE_LUT_2936 16'h2935
`define CUBE_LUT_2937 16'h2936
`define CUBE_LUT_2938 16'h2937
`define CUBE_LUT_2939 16'h2938
`define CUBE_LUT_293A 16'h2939
`define CUBE_LUT_293B 16'h293A
`define CUBE_LUT_293C 16'h293B
`define CUBE_LUT_293D 16'h293C
`define CUBE_LUT_293E 16'h293D
`define CUBE_LUT_293F 16'h293E
`define CUBE_LUT_2940 16'h293F
`define CUBE_LUT_2941 16'h2940
`define CUBE_LUT_2942 16'h2941
`define CUBE_LUT_2943 16'h2942
`define CUBE_LUT_2944 16'h2943
`define CUBE_LUT_2945 16'h2944
`define CUBE_LUT_2946 16'h2945
`define CUBE_LUT_2947 16'h2946
`define CUBE_LUT_2948 16'h2947
`define CUBE_LUT_2949 16'h2948
`define CUBE_LUT_294A 16'h2949
`define CUBE_LUT_294B 16'h294A
`define CUBE_LUT_294C 16'h294B
`define CUBE_LUT_294D 16'h294C
`define CUBE_LUT_294E 16'h294D
`define CUBE_LUT_294F 16'h294E
`define CUBE_LUT_2950 16'h294F
`define CUBE_LUT_2951 16'h2950
`define CUBE_LUT_2952 16'h2951
`define CUBE_LUT_2953 16'h2952
`define CUBE_LUT_2954 16'h2953
`define CUBE_LUT_2955 16'h2954
`define CUBE_LUT_2956 16'h2955
`define CUBE_LUT_2957 16'h2956
`define CUBE_LUT_2958 16'h2957
`define CUBE_LUT_2959 16'h2958
`define CUBE_LUT_295A 16'h2959
`define CUBE_LUT_295B 16'h295A
`define CUBE_LUT_295C 16'h295B
`define CUBE_LUT_295D 16'h295C
`define CUBE_LUT_295E 16'h295D
`define CUBE_LUT_295F 16'h295E
`define CUBE_LUT_2960 16'h295F
`define CUBE_LUT_2961 16'h2960
`define CUBE_LUT_2962 16'h2961
`define CUBE_LUT_2963 16'h2962
`define CUBE_LUT_2964 16'h2963
`define CUBE_LUT_2965 16'h2964
`define CUBE_LUT_2966 16'h2965
`define CUBE_LUT_2967 16'h2966
`define CUBE_LUT_2968 16'h2967
`define CUBE_LUT_2969 16'h2968
`define CUBE_LUT_296A 16'h2969
`define CUBE_LUT_296B 16'h296A
`define CUBE_LUT_296C 16'h296B
`define CUBE_LUT_296D 16'h296C
`define CUBE_LUT_296E 16'h296D
`define CUBE_LUT_296F 16'h296E
`define CUBE_LUT_2970 16'h296F
`define CUBE_LUT_2971 16'h2970
`define CUBE_LUT_2972 16'h2971
`define CUBE_LUT_2973 16'h2972
`define CUBE_LUT_2974 16'h2973
`define CUBE_LUT_2975 16'h2974
`define CUBE_LUT_2976 16'h2975
`define CUBE_LUT_2977 16'h2976
`define CUBE_LUT_2978 16'h2977
`define CUBE_LUT_2979 16'h2978
`define CUBE_LUT_297A 16'h2979
`define CUBE_LUT_297B 16'h297A
`define CUBE_LUT_297C 16'h297B
`define CUBE_LUT_297D 16'h297C
`define CUBE_LUT_297E 16'h297D
`define CUBE_LUT_297F 16'h297E
`define CUBE_LUT_2980 16'h297F
`define CUBE_LUT_2981 16'h2980
`define CUBE_LUT_2982 16'h2981
`define CUBE_LUT_2983 16'h2982
`define CUBE_LUT_2984 16'h2983
`define CUBE_LUT_2985 16'h2984
`define CUBE_LUT_2986 16'h2985
`define CUBE_LUT_2987 16'h2986
`define CUBE_LUT_2988 16'h2987
`define CUBE_LUT_2989 16'h2988
`define CUBE_LUT_298A 16'h2989
`define CUBE_LUT_298B 16'h298A
`define CUBE_LUT_298C 16'h298B
`define CUBE_LUT_298D 16'h298C
`define CUBE_LUT_298E 16'h298D
`define CUBE_LUT_298F 16'h298E
`define CUBE_LUT_2990 16'h298F
`define CUBE_LUT_2991 16'h2990
`define CUBE_LUT_2992 16'h2991
`define CUBE_LUT_2993 16'h2992
`define CUBE_LUT_2994 16'h2993
`define CUBE_LUT_2995 16'h2994
`define CUBE_LUT_2996 16'h2995
`define CUBE_LUT_2997 16'h2996
`define CUBE_LUT_2998 16'h2997
`define CUBE_LUT_2999 16'h2998
`define CUBE_LUT_299A 16'h2999
`define CUBE_LUT_299B 16'h299A
`define CUBE_LUT_299C 16'h299B
`define CUBE_LUT_299D 16'h299C
`define CUBE_LUT_299E 16'h299D
`define CUBE_LUT_299F 16'h299E
`define CUBE_LUT_29A0 16'h299F
`define CUBE_LUT_29A1 16'h29A0
`define CUBE_LUT_29A2 16'h29A1
`define CUBE_LUT_29A3 16'h29A2
`define CUBE_LUT_29A4 16'h29A3
`define CUBE_LUT_29A5 16'h29A4
`define CUBE_LUT_29A6 16'h29A5
`define CUBE_LUT_29A7 16'h29A6
`define CUBE_LUT_29A8 16'h29A7
`define CUBE_LUT_29A9 16'h29A8
`define CUBE_LUT_29AA 16'h29A9
`define CUBE_LUT_29AB 16'h29AA
`define CUBE_LUT_29AC 16'h29AB
`define CUBE_LUT_29AD 16'h29AC
`define CUBE_LUT_29AE 16'h29AD
`define CUBE_LUT_29AF 16'h29AE
`define CUBE_LUT_29B0 16'h29AF
`define CUBE_LUT_29B1 16'h29B0
`define CUBE_LUT_29B2 16'h29B1
`define CUBE_LUT_29B3 16'h29B2
`define CUBE_LUT_29B4 16'h29B3
`define CUBE_LUT_29B5 16'h29B4
`define CUBE_LUT_29B6 16'h29B5
`define CUBE_LUT_29B7 16'h29B6
`define CUBE_LUT_29B8 16'h29B7
`define CUBE_LUT_29B9 16'h29B8
`define CUBE_LUT_29BA 16'h29B9
`define CUBE_LUT_29BB 16'h29BA
`define CUBE_LUT_29BC 16'h29BB
`define CUBE_LUT_29BD 16'h29BC
`define CUBE_LUT_29BE 16'h29BD
`define CUBE_LUT_29BF 16'h29BE
`define CUBE_LUT_29C0 16'h29BF
`define CUBE_LUT_29C1 16'h29C0
`define CUBE_LUT_29C2 16'h29C1
`define CUBE_LUT_29C3 16'h29C2
`define CUBE_LUT_29C4 16'h29C3
`define CUBE_LUT_29C5 16'h29C4
`define CUBE_LUT_29C6 16'h29C5
`define CUBE_LUT_29C7 16'h29C6
`define CUBE_LUT_29C8 16'h29C7
`define CUBE_LUT_29C9 16'h29C8
`define CUBE_LUT_29CA 16'h29C9
`define CUBE_LUT_29CB 16'h29CA
`define CUBE_LUT_29CC 16'h29CB
`define CUBE_LUT_29CD 16'h29CC
`define CUBE_LUT_29CE 16'h29CD
`define CUBE_LUT_29CF 16'h29CE
`define CUBE_LUT_29D0 16'h29CF
`define CUBE_LUT_29D1 16'h29D0
`define CUBE_LUT_29D2 16'h29D1
`define CUBE_LUT_29D3 16'h29D2
`define CUBE_LUT_29D4 16'h29D3
`define CUBE_LUT_29D5 16'h29D4
`define CUBE_LUT_29D6 16'h29D5
`define CUBE_LUT_29D7 16'h29D6
`define CUBE_LUT_29D8 16'h29D7
`define CUBE_LUT_29D9 16'h29D8
`define CUBE_LUT_29DA 16'h29D9
`define CUBE_LUT_29DB 16'h29DA
`define CUBE_LUT_29DC 16'h29DB
`define CUBE_LUT_29DD 16'h29DC
`define CUBE_LUT_29DE 16'h29DD
`define CUBE_LUT_29DF 16'h29DE
`define CUBE_LUT_29E0 16'h29DF
`define CUBE_LUT_29E1 16'h29E0
`define CUBE_LUT_29E2 16'h29E1
`define CUBE_LUT_29E3 16'h29E2
`define CUBE_LUT_29E4 16'h29E3
`define CUBE_LUT_29E5 16'h29E4
`define CUBE_LUT_29E6 16'h29E5
`define CUBE_LUT_29E7 16'h29E6
`define CUBE_LUT_29E8 16'h29E7
`define CUBE_LUT_29E9 16'h29E8
`define CUBE_LUT_29EA 16'h29E9
`define CUBE_LUT_29EB 16'h29EA
`define CUBE_LUT_29EC 16'h29EB
`define CUBE_LUT_29ED 16'h29EC
`define CUBE_LUT_29EE 16'h29ED
`define CUBE_LUT_29EF 16'h29EE
`define CUBE_LUT_29F0 16'h29EF
`define CUBE_LUT_29F1 16'h29F0
`define CUBE_LUT_29F2 16'h29F1
`define CUBE_LUT_29F3 16'h29F2
`define CUBE_LUT_29F4 16'h29F3
`define CUBE_LUT_29F5 16'h29F4
`define CUBE_LUT_29F6 16'h29F5
`define CUBE_LUT_29F7 16'h29F6
`define CUBE_LUT_29F8 16'h29F7
`define CUBE_LUT_29F9 16'h29F8
`define CUBE_LUT_29FA 16'h29F9
`define CUBE_LUT_29FB 16'h29FA
`define CUBE_LUT_29FC 16'h29FB
`define CUBE_LUT_29FD 16'h29FC
`define CUBE_LUT_29FE 16'h29FD
`define CUBE_LUT_29FF 16'h29FE
`define CUBE_LUT_2A00 16'h29FF
`define CUBE_LUT_2A01 16'h2A00
`define CUBE_LUT_2A02 16'h2A01
`define CUBE_LUT_2A03 16'h2A02
`define CUBE_LUT_2A04 16'h2A03
`define CUBE_LUT_2A05 16'h2A04
`define CUBE_LUT_2A06 16'h2A05
`define CUBE_LUT_2A07 16'h2A06
`define CUBE_LUT_2A08 16'h2A07
`define CUBE_LUT_2A09 16'h2A08
`define CUBE_LUT_2A0A 16'h2A09
`define CUBE_LUT_2A0B 16'h2A0A
`define CUBE_LUT_2A0C 16'h2A0B
`define CUBE_LUT_2A0D 16'h2A0C
`define CUBE_LUT_2A0E 16'h2A0D
`define CUBE_LUT_2A0F 16'h2A0E
`define CUBE_LUT_2A10 16'h2A0F
`define CUBE_LUT_2A11 16'h2A10
`define CUBE_LUT_2A12 16'h2A11
`define CUBE_LUT_2A13 16'h2A12
`define CUBE_LUT_2A14 16'h2A13
`define CUBE_LUT_2A15 16'h2A14
`define CUBE_LUT_2A16 16'h2A15
`define CUBE_LUT_2A17 16'h2A16
`define CUBE_LUT_2A18 16'h2A17
`define CUBE_LUT_2A19 16'h2A18
`define CUBE_LUT_2A1A 16'h2A19
`define CUBE_LUT_2A1B 16'h2A1A
`define CUBE_LUT_2A1C 16'h2A1B
`define CUBE_LUT_2A1D 16'h2A1C
`define CUBE_LUT_2A1E 16'h2A1D
`define CUBE_LUT_2A1F 16'h2A1E
`define CUBE_LUT_2A20 16'h2A1F
`define CUBE_LUT_2A21 16'h2A20
`define CUBE_LUT_2A22 16'h2A21
`define CUBE_LUT_2A23 16'h2A22
`define CUBE_LUT_2A24 16'h2A23
`define CUBE_LUT_2A25 16'h2A24
`define CUBE_LUT_2A26 16'h2A25
`define CUBE_LUT_2A27 16'h2A26
`define CUBE_LUT_2A28 16'h2A27
`define CUBE_LUT_2A29 16'h2A28
`define CUBE_LUT_2A2A 16'h2A29
`define CUBE_LUT_2A2B 16'h2A2A
`define CUBE_LUT_2A2C 16'h2A2B
`define CUBE_LUT_2A2D 16'h2A2C
`define CUBE_LUT_2A2E 16'h2A2D
`define CUBE_LUT_2A2F 16'h2A2E
`define CUBE_LUT_2A30 16'h2A2F
`define CUBE_LUT_2A31 16'h2A30
`define CUBE_LUT_2A32 16'h2A31
`define CUBE_LUT_2A33 16'h2A32
`define CUBE_LUT_2A34 16'h2A33
`define CUBE_LUT_2A35 16'h2A34
`define CUBE_LUT_2A36 16'h2A35
`define CUBE_LUT_2A37 16'h2A36
`define CUBE_LUT_2A38 16'h2A37
`define CUBE_LUT_2A39 16'h2A38
`define CUBE_LUT_2A3A 16'h2A39
`define CUBE_LUT_2A3B 16'h2A3A
`define CUBE_LUT_2A3C 16'h2A3B
`define CUBE_LUT_2A3D 16'h2A3C
`define CUBE_LUT_2A3E 16'h2A3D
`define CUBE_LUT_2A3F 16'h2A3E
`define CUBE_LUT_2A40 16'h2A3F
`define CUBE_LUT_2A41 16'h2A40
`define CUBE_LUT_2A42 16'h2A41
`define CUBE_LUT_2A43 16'h2A42
`define CUBE_LUT_2A44 16'h2A43
`define CUBE_LUT_2A45 16'h2A44
`define CUBE_LUT_2A46 16'h2A45
`define CUBE_LUT_2A47 16'h2A46
`define CUBE_LUT_2A48 16'h2A47
`define CUBE_LUT_2A49 16'h2A48
`define CUBE_LUT_2A4A 16'h2A49
`define CUBE_LUT_2A4B 16'h2A4A
`define CUBE_LUT_2A4C 16'h2A4B
`define CUBE_LUT_2A4D 16'h2A4C
`define CUBE_LUT_2A4E 16'h2A4D
`define CUBE_LUT_2A4F 16'h2A4E
`define CUBE_LUT_2A50 16'h2A4F
`define CUBE_LUT_2A51 16'h2A50
`define CUBE_LUT_2A52 16'h2A51
`define CUBE_LUT_2A53 16'h2A52
`define CUBE_LUT_2A54 16'h2A53
`define CUBE_LUT_2A55 16'h2A54
`define CUBE_LUT_2A56 16'h2A55
`define CUBE_LUT_2A57 16'h2A56
`define CUBE_LUT_2A58 16'h2A57
`define CUBE_LUT_2A59 16'h2A58
`define CUBE_LUT_2A5A 16'h2A59
`define CUBE_LUT_2A5B 16'h2A5A
`define CUBE_LUT_2A5C 16'h2A5B
`define CUBE_LUT_2A5D 16'h2A5C
`define CUBE_LUT_2A5E 16'h2A5D
`define CUBE_LUT_2A5F 16'h2A5E
`define CUBE_LUT_2A60 16'h2A5F
`define CUBE_LUT_2A61 16'h2A60
`define CUBE_LUT_2A62 16'h2A61
`define CUBE_LUT_2A63 16'h2A62
`define CUBE_LUT_2A64 16'h2A63
`define CUBE_LUT_2A65 16'h2A64
`define CUBE_LUT_2A66 16'h2A65
`define CUBE_LUT_2A67 16'h2A66
`define CUBE_LUT_2A68 16'h2A67
`define CUBE_LUT_2A69 16'h2A68
`define CUBE_LUT_2A6A 16'h2A69
`define CUBE_LUT_2A6B 16'h2A6A
`define CUBE_LUT_2A6C 16'h2A6B
`define CUBE_LUT_2A6D 16'h2A6C
`define CUBE_LUT_2A6E 16'h2A6D
`define CUBE_LUT_2A6F 16'h2A6E
`define CUBE_LUT_2A70 16'h2A6F
`define CUBE_LUT_2A71 16'h2A70
`define CUBE_LUT_2A72 16'h2A71
`define CUBE_LUT_2A73 16'h2A72
`define CUBE_LUT_2A74 16'h2A73
`define CUBE_LUT_2A75 16'h2A74
`define CUBE_LUT_2A76 16'h2A75
`define CUBE_LUT_2A77 16'h2A76
`define CUBE_LUT_2A78 16'h2A77
`define CUBE_LUT_2A79 16'h2A78
`define CUBE_LUT_2A7A 16'h2A79
`define CUBE_LUT_2A7B 16'h2A7A
`define CUBE_LUT_2A7C 16'h2A7B
`define CUBE_LUT_2A7D 16'h2A7C
`define CUBE_LUT_2A7E 16'h2A7D
`define CUBE_LUT_2A7F 16'h2A7E
`define CUBE_LUT_2A80 16'h2A7F
`define CUBE_LUT_2A81 16'h2A80
`define CUBE_LUT_2A82 16'h2A81
`define CUBE_LUT_2A83 16'h2A82
`define CUBE_LUT_2A84 16'h2A83
`define CUBE_LUT_2A85 16'h2A84
`define CUBE_LUT_2A86 16'h2A85
`define CUBE_LUT_2A87 16'h2A86
`define CUBE_LUT_2A88 16'h2A87
`define CUBE_LUT_2A89 16'h2A88
`define CUBE_LUT_2A8A 16'h2A89
`define CUBE_LUT_2A8B 16'h2A8A
`define CUBE_LUT_2A8C 16'h2A8B
`define CUBE_LUT_2A8D 16'h2A8C
`define CUBE_LUT_2A8E 16'h2A8D
`define CUBE_LUT_2A8F 16'h2A8E
`define CUBE_LUT_2A90 16'h2A8F
`define CUBE_LUT_2A91 16'h2A90
`define CUBE_LUT_2A92 16'h2A91
`define CUBE_LUT_2A93 16'h2A92
`define CUBE_LUT_2A94 16'h2A93
`define CUBE_LUT_2A95 16'h2A94
`define CUBE_LUT_2A96 16'h2A95
`define CUBE_LUT_2A97 16'h2A96
`define CUBE_LUT_2A98 16'h2A97
`define CUBE_LUT_2A99 16'h2A98
`define CUBE_LUT_2A9A 16'h2A99
`define CUBE_LUT_2A9B 16'h2A9A
`define CUBE_LUT_2A9C 16'h2A9A
`define CUBE_LUT_2A9D 16'h2A9B
`define CUBE_LUT_2A9E 16'h2A9C
`define CUBE_LUT_2A9F 16'h2A9D
`define CUBE_LUT_2AA0 16'h2A9E
`define CUBE_LUT_2AA1 16'h2A9F
`define CUBE_LUT_2AA2 16'h2AA0
`define CUBE_LUT_2AA3 16'h2AA1
`define CUBE_LUT_2AA4 16'h2AA2
`define CUBE_LUT_2AA5 16'h2AA3
`define CUBE_LUT_2AA6 16'h2AA4
`define CUBE_LUT_2AA7 16'h2AA5
`define CUBE_LUT_2AA8 16'h2AA6
`define CUBE_LUT_2AA9 16'h2AA7
`define CUBE_LUT_2AAA 16'h2AA8
`define CUBE_LUT_2AAB 16'h2AA9
`define CUBE_LUT_2AAC 16'h2AAA
`define CUBE_LUT_2AAD 16'h2AAB
`define CUBE_LUT_2AAE 16'h2AAC
`define CUBE_LUT_2AAF 16'h2AAD
`define CUBE_LUT_2AB0 16'h2AAE
`define CUBE_LUT_2AB1 16'h2AAF
`define CUBE_LUT_2AB2 16'h2AB0
`define CUBE_LUT_2AB3 16'h2AB1
`define CUBE_LUT_2AB4 16'h2AB2
`define CUBE_LUT_2AB5 16'h2AB3
`define CUBE_LUT_2AB6 16'h2AB4
`define CUBE_LUT_2AB7 16'h2AB5
`define CUBE_LUT_2AB8 16'h2AB6
`define CUBE_LUT_2AB9 16'h2AB7
`define CUBE_LUT_2ABA 16'h2AB8
`define CUBE_LUT_2ABB 16'h2AB9
`define CUBE_LUT_2ABC 16'h2ABA
`define CUBE_LUT_2ABD 16'h2ABB
`define CUBE_LUT_2ABE 16'h2ABC
`define CUBE_LUT_2ABF 16'h2ABD
`define CUBE_LUT_2AC0 16'h2ABE
`define CUBE_LUT_2AC1 16'h2ABF
`define CUBE_LUT_2AC2 16'h2AC0
`define CUBE_LUT_2AC3 16'h2AC1
`define CUBE_LUT_2AC4 16'h2AC2
`define CUBE_LUT_2AC5 16'h2AC3
`define CUBE_LUT_2AC6 16'h2AC4
`define CUBE_LUT_2AC7 16'h2AC5
`define CUBE_LUT_2AC8 16'h2AC6
`define CUBE_LUT_2AC9 16'h2AC7
`define CUBE_LUT_2ACA 16'h2AC8
`define CUBE_LUT_2ACB 16'h2AC9
`define CUBE_LUT_2ACC 16'h2ACA
`define CUBE_LUT_2ACD 16'h2ACB
`define CUBE_LUT_2ACE 16'h2ACC
`define CUBE_LUT_2ACF 16'h2ACD
`define CUBE_LUT_2AD0 16'h2ACE
`define CUBE_LUT_2AD1 16'h2ACF
`define CUBE_LUT_2AD2 16'h2AD0
`define CUBE_LUT_2AD3 16'h2AD1
`define CUBE_LUT_2AD4 16'h2AD2
`define CUBE_LUT_2AD5 16'h2AD3
`define CUBE_LUT_2AD6 16'h2AD4
`define CUBE_LUT_2AD7 16'h2AD5
`define CUBE_LUT_2AD8 16'h2AD6
`define CUBE_LUT_2AD9 16'h2AD7
`define CUBE_LUT_2ADA 16'h2AD8
`define CUBE_LUT_2ADB 16'h2AD9
`define CUBE_LUT_2ADC 16'h2ADA
`define CUBE_LUT_2ADD 16'h2ADB
`define CUBE_LUT_2ADE 16'h2ADC
`define CUBE_LUT_2ADF 16'h2ADD
`define CUBE_LUT_2AE0 16'h2ADE
`define CUBE_LUT_2AE1 16'h2ADF
`define CUBE_LUT_2AE2 16'h2AE0
`define CUBE_LUT_2AE3 16'h2AE1
`define CUBE_LUT_2AE4 16'h2AE2
`define CUBE_LUT_2AE5 16'h2AE3
`define CUBE_LUT_2AE6 16'h2AE4
`define CUBE_LUT_2AE7 16'h2AE5
`define CUBE_LUT_2AE8 16'h2AE6
`define CUBE_LUT_2AE9 16'h2AE7
`define CUBE_LUT_2AEA 16'h2AE8
`define CUBE_LUT_2AEB 16'h2AE9
`define CUBE_LUT_2AEC 16'h2AEA
`define CUBE_LUT_2AED 16'h2AEB
`define CUBE_LUT_2AEE 16'h2AEC
`define CUBE_LUT_2AEF 16'h2AED
`define CUBE_LUT_2AF0 16'h2AEE
`define CUBE_LUT_2AF1 16'h2AEF
`define CUBE_LUT_2AF2 16'h2AF0
`define CUBE_LUT_2AF3 16'h2AF1
`define CUBE_LUT_2AF4 16'h2AF2
`define CUBE_LUT_2AF5 16'h2AF3
`define CUBE_LUT_2AF6 16'h2AF4
`define CUBE_LUT_2AF7 16'h2AF5
`define CUBE_LUT_2AF8 16'h2AF6
`define CUBE_LUT_2AF9 16'h2AF7
`define CUBE_LUT_2AFA 16'h2AF8
`define CUBE_LUT_2AFB 16'h2AF9
`define CUBE_LUT_2AFC 16'h2AFA
`define CUBE_LUT_2AFD 16'h2AFB
`define CUBE_LUT_2AFE 16'h2AFC
`define CUBE_LUT_2AFF 16'h2AFD
`define CUBE_LUT_2B00 16'h2AFE
`define CUBE_LUT_2B01 16'h2AFF
`define CUBE_LUT_2B02 16'h2B00
`define CUBE_LUT_2B03 16'h2B01
`define CUBE_LUT_2B04 16'h2B02
`define CUBE_LUT_2B05 16'h2B03
`define CUBE_LUT_2B06 16'h2B04
`define CUBE_LUT_2B07 16'h2B05
`define CUBE_LUT_2B08 16'h2B06
`define CUBE_LUT_2B09 16'h2B07
`define CUBE_LUT_2B0A 16'h2B08
`define CUBE_LUT_2B0B 16'h2B09
`define CUBE_LUT_2B0C 16'h2B0A
`define CUBE_LUT_2B0D 16'h2B0B
`define CUBE_LUT_2B0E 16'h2B0C
`define CUBE_LUT_2B0F 16'h2B0D
`define CUBE_LUT_2B10 16'h2B0E
`define CUBE_LUT_2B11 16'h2B0F
`define CUBE_LUT_2B12 16'h2B10
`define CUBE_LUT_2B13 16'h2B11
`define CUBE_LUT_2B14 16'h2B12
`define CUBE_LUT_2B15 16'h2B13
`define CUBE_LUT_2B16 16'h2B14
`define CUBE_LUT_2B17 16'h2B15
`define CUBE_LUT_2B18 16'h2B16
`define CUBE_LUT_2B19 16'h2B17
`define CUBE_LUT_2B1A 16'h2B18
`define CUBE_LUT_2B1B 16'h2B19
`define CUBE_LUT_2B1C 16'h2B1A
`define CUBE_LUT_2B1D 16'h2B1B
`define CUBE_LUT_2B1E 16'h2B1C
`define CUBE_LUT_2B1F 16'h2B1D
`define CUBE_LUT_2B20 16'h2B1E
`define CUBE_LUT_2B21 16'h2B1F
`define CUBE_LUT_2B22 16'h2B20
`define CUBE_LUT_2B23 16'h2B21
`define CUBE_LUT_2B24 16'h2B22
`define CUBE_LUT_2B25 16'h2B23
`define CUBE_LUT_2B26 16'h2B24
`define CUBE_LUT_2B27 16'h2B25
`define CUBE_LUT_2B28 16'h2B26
`define CUBE_LUT_2B29 16'h2B27
`define CUBE_LUT_2B2A 16'h2B28
`define CUBE_LUT_2B2B 16'h2B29
`define CUBE_LUT_2B2C 16'h2B2A
`define CUBE_LUT_2B2D 16'h2B2B
`define CUBE_LUT_2B2E 16'h2B2C
`define CUBE_LUT_2B2F 16'h2B2D
`define CUBE_LUT_2B30 16'h2B2E
`define CUBE_LUT_2B31 16'h2B2F
`define CUBE_LUT_2B32 16'h2B30
`define CUBE_LUT_2B33 16'h2B31
`define CUBE_LUT_2B34 16'h2B32
`define CUBE_LUT_2B35 16'h2B33
`define CUBE_LUT_2B36 16'h2B34
`define CUBE_LUT_2B37 16'h2B35
`define CUBE_LUT_2B38 16'h2B36
`define CUBE_LUT_2B39 16'h2B37
`define CUBE_LUT_2B3A 16'h2B38
`define CUBE_LUT_2B3B 16'h2B39
`define CUBE_LUT_2B3C 16'h2B3A
`define CUBE_LUT_2B3D 16'h2B3B
`define CUBE_LUT_2B3E 16'h2B3C
`define CUBE_LUT_2B3F 16'h2B3D
`define CUBE_LUT_2B40 16'h2B3E
`define CUBE_LUT_2B41 16'h2B3F
`define CUBE_LUT_2B42 16'h2B40
`define CUBE_LUT_2B43 16'h2B41
`define CUBE_LUT_2B44 16'h2B42
`define CUBE_LUT_2B45 16'h2B43
`define CUBE_LUT_2B46 16'h2B44
`define CUBE_LUT_2B47 16'h2B45
`define CUBE_LUT_2B48 16'h2B46
`define CUBE_LUT_2B49 16'h2B47
`define CUBE_LUT_2B4A 16'h2B48
`define CUBE_LUT_2B4B 16'h2B49
`define CUBE_LUT_2B4C 16'h2B4A
`define CUBE_LUT_2B4D 16'h2B4B
`define CUBE_LUT_2B4E 16'h2B4C
`define CUBE_LUT_2B4F 16'h2B4D
`define CUBE_LUT_2B50 16'h2B4E
`define CUBE_LUT_2B51 16'h2B4F
`define CUBE_LUT_2B52 16'h2B50
`define CUBE_LUT_2B53 16'h2B51
`define CUBE_LUT_2B54 16'h2B52
`define CUBE_LUT_2B55 16'h2B53
`define CUBE_LUT_2B56 16'h2B54
`define CUBE_LUT_2B57 16'h2B55
`define CUBE_LUT_2B58 16'h2B56
`define CUBE_LUT_2B59 16'h2B57
`define CUBE_LUT_2B5A 16'h2B58
`define CUBE_LUT_2B5B 16'h2B59
`define CUBE_LUT_2B5C 16'h2B5A
`define CUBE_LUT_2B5D 16'h2B5B
`define CUBE_LUT_2B5E 16'h2B5C
`define CUBE_LUT_2B5F 16'h2B5D
`define CUBE_LUT_2B60 16'h2B5E
`define CUBE_LUT_2B61 16'h2B5F
`define CUBE_LUT_2B62 16'h2B60
`define CUBE_LUT_2B63 16'h2B61
`define CUBE_LUT_2B64 16'h2B62
`define CUBE_LUT_2B65 16'h2B63
`define CUBE_LUT_2B66 16'h2B64
`define CUBE_LUT_2B67 16'h2B65
`define CUBE_LUT_2B68 16'h2B66
`define CUBE_LUT_2B69 16'h2B67
`define CUBE_LUT_2B6A 16'h2B68
`define CUBE_LUT_2B6B 16'h2B69
`define CUBE_LUT_2B6C 16'h2B6A
`define CUBE_LUT_2B6D 16'h2B6B
`define CUBE_LUT_2B6E 16'h2B6C
`define CUBE_LUT_2B6F 16'h2B6D
`define CUBE_LUT_2B70 16'h2B6E
`define CUBE_LUT_2B71 16'h2B6F
`define CUBE_LUT_2B72 16'h2B70
`define CUBE_LUT_2B73 16'h2B71
`define CUBE_LUT_2B74 16'h2B72
`define CUBE_LUT_2B75 16'h2B73
`define CUBE_LUT_2B76 16'h2B74
`define CUBE_LUT_2B77 16'h2B75
`define CUBE_LUT_2B78 16'h2B76
`define CUBE_LUT_2B79 16'h2B77
`define CUBE_LUT_2B7A 16'h2B78
`define CUBE_LUT_2B7B 16'h2B79
`define CUBE_LUT_2B7C 16'h2B7A
`define CUBE_LUT_2B7D 16'h2B7B
`define CUBE_LUT_2B7E 16'h2B7C
`define CUBE_LUT_2B7F 16'h2B7D
`define CUBE_LUT_2B80 16'h2B7E
`define CUBE_LUT_2B81 16'h2B7F
`define CUBE_LUT_2B82 16'h2B80
`define CUBE_LUT_2B83 16'h2B81
`define CUBE_LUT_2B84 16'h2B82
`define CUBE_LUT_2B85 16'h2B83
`define CUBE_LUT_2B86 16'h2B84
`define CUBE_LUT_2B87 16'h2B85
`define CUBE_LUT_2B88 16'h2B86
`define CUBE_LUT_2B89 16'h2B87
`define CUBE_LUT_2B8A 16'h2B88
`define CUBE_LUT_2B8B 16'h2B89
`define CUBE_LUT_2B8C 16'h2B8A
`define CUBE_LUT_2B8D 16'h2B8B
`define CUBE_LUT_2B8E 16'h2B8C
`define CUBE_LUT_2B8F 16'h2B8D
`define CUBE_LUT_2B90 16'h2B8E
`define CUBE_LUT_2B91 16'h2B8F
`define CUBE_LUT_2B92 16'h2B90
`define CUBE_LUT_2B93 16'h2B91
`define CUBE_LUT_2B94 16'h2B92
`define CUBE_LUT_2B95 16'h2B93
`define CUBE_LUT_2B96 16'h2B94
`define CUBE_LUT_2B97 16'h2B95
`define CUBE_LUT_2B98 16'h2B96
`define CUBE_LUT_2B99 16'h2B97
`define CUBE_LUT_2B9A 16'h2B98
`define CUBE_LUT_2B9B 16'h2B99
`define CUBE_LUT_2B9C 16'h2B9A
`define CUBE_LUT_2B9D 16'h2B9B
`define CUBE_LUT_2B9E 16'h2B9C
`define CUBE_LUT_2B9F 16'h2B9D
`define CUBE_LUT_2BA0 16'h2B9E
`define CUBE_LUT_2BA1 16'h2B9F
`define CUBE_LUT_2BA2 16'h2BA0
`define CUBE_LUT_2BA3 16'h2BA1
`define CUBE_LUT_2BA4 16'h2BA2
`define CUBE_LUT_2BA5 16'h2BA3
`define CUBE_LUT_2BA6 16'h2BA4
`define CUBE_LUT_2BA7 16'h2BA5
`define CUBE_LUT_2BA8 16'h2BA6
`define CUBE_LUT_2BA9 16'h2BA7
`define CUBE_LUT_2BAA 16'h2BA8
`define CUBE_LUT_2BAB 16'h2BA9
`define CUBE_LUT_2BAC 16'h2BAA
`define CUBE_LUT_2BAD 16'h2BAB
`define CUBE_LUT_2BAE 16'h2BAC
`define CUBE_LUT_2BAF 16'h2BAD
`define CUBE_LUT_2BB0 16'h2BAE
`define CUBE_LUT_2BB1 16'h2BAF
`define CUBE_LUT_2BB2 16'h2BB0
`define CUBE_LUT_2BB3 16'h2BB1
`define CUBE_LUT_2BB4 16'h2BB2
`define CUBE_LUT_2BB5 16'h2BB3
`define CUBE_LUT_2BB6 16'h2BB4
`define CUBE_LUT_2BB7 16'h2BB5
`define CUBE_LUT_2BB8 16'h2BB6
`define CUBE_LUT_2BB9 16'h2BB7
`define CUBE_LUT_2BBA 16'h2BB8
`define CUBE_LUT_2BBB 16'h2BB9
`define CUBE_LUT_2BBC 16'h2BBA
`define CUBE_LUT_2BBD 16'h2BBB
`define CUBE_LUT_2BBE 16'h2BBC
`define CUBE_LUT_2BBF 16'h2BBD
`define CUBE_LUT_2BC0 16'h2BBE
`define CUBE_LUT_2BC1 16'h2BBF
`define CUBE_LUT_2BC2 16'h2BC0
`define CUBE_LUT_2BC3 16'h2BC1
`define CUBE_LUT_2BC4 16'h2BC2
`define CUBE_LUT_2BC5 16'h2BC3
`define CUBE_LUT_2BC6 16'h2BC4
`define CUBE_LUT_2BC7 16'h2BC5
`define CUBE_LUT_2BC8 16'h2BC6
`define CUBE_LUT_2BC9 16'h2BC7
`define CUBE_LUT_2BCA 16'h2BC8
`define CUBE_LUT_2BCB 16'h2BC9
`define CUBE_LUT_2BCC 16'h2BCA
`define CUBE_LUT_2BCD 16'h2BCB
`define CUBE_LUT_2BCE 16'h2BCC
`define CUBE_LUT_2BCF 16'h2BCD
`define CUBE_LUT_2BD0 16'h2BCE
`define CUBE_LUT_2BD1 16'h2BCF
`define CUBE_LUT_2BD2 16'h2BD0
`define CUBE_LUT_2BD3 16'h2BD1
`define CUBE_LUT_2BD4 16'h2BD2
`define CUBE_LUT_2BD5 16'h2BD3
`define CUBE_LUT_2BD6 16'h2BD3
`define CUBE_LUT_2BD7 16'h2BD4
`define CUBE_LUT_2BD8 16'h2BD5
`define CUBE_LUT_2BD9 16'h2BD6
`define CUBE_LUT_2BDA 16'h2BD7
`define CUBE_LUT_2BDB 16'h2BD8
`define CUBE_LUT_2BDC 16'h2BD9
`define CUBE_LUT_2BDD 16'h2BDA
`define CUBE_LUT_2BDE 16'h2BDB
`define CUBE_LUT_2BDF 16'h2BDC
`define CUBE_LUT_2BE0 16'h2BDD
`define CUBE_LUT_2BE1 16'h2BDE
`define CUBE_LUT_2BE2 16'h2BDF
`define CUBE_LUT_2BE3 16'h2BE0
`define CUBE_LUT_2BE4 16'h2BE1
`define CUBE_LUT_2BE5 16'h2BE2
`define CUBE_LUT_2BE6 16'h2BE3
`define CUBE_LUT_2BE7 16'h2BE4
`define CUBE_LUT_2BE8 16'h2BE5
`define CUBE_LUT_2BE9 16'h2BE6
`define CUBE_LUT_2BEA 16'h2BE7
`define CUBE_LUT_2BEB 16'h2BE8
`define CUBE_LUT_2BEC 16'h2BE9
`define CUBE_LUT_2BED 16'h2BEA
`define CUBE_LUT_2BEE 16'h2BEB
`define CUBE_LUT_2BEF 16'h2BEC
`define CUBE_LUT_2BF0 16'h2BED
`define CUBE_LUT_2BF1 16'h2BEE
`define CUBE_LUT_2BF2 16'h2BEF
`define CUBE_LUT_2BF3 16'h2BF0
`define CUBE_LUT_2BF4 16'h2BF1
`define CUBE_LUT_2BF5 16'h2BF2
`define CUBE_LUT_2BF6 16'h2BF3
`define CUBE_LUT_2BF7 16'h2BF4
`define CUBE_LUT_2BF8 16'h2BF5
`define CUBE_LUT_2BF9 16'h2BF6
`define CUBE_LUT_2BFA 16'h2BF7
`define CUBE_LUT_2BFB 16'h2BF8
`define CUBE_LUT_2BFC 16'h2BF9
`define CUBE_LUT_2BFD 16'h2BFA
`define CUBE_LUT_2BFE 16'h2BFB
`define CUBE_LUT_2BFF 16'h2BFC
`define CUBE_LUT_2C00 16'h2BFD
`define CUBE_LUT_2C01 16'h2BFF
`define CUBE_LUT_2C02 16'h2C01
`define CUBE_LUT_2C03 16'h2C02
`define CUBE_LUT_2C04 16'h2C03
`define CUBE_LUT_2C05 16'h2C04
`define CUBE_LUT_2C06 16'h2C05
`define CUBE_LUT_2C07 16'h2C06
`define CUBE_LUT_2C08 16'h2C07
`define CUBE_LUT_2C09 16'h2C08
`define CUBE_LUT_2C0A 16'h2C09
`define CUBE_LUT_2C0B 16'h2C0A
`define CUBE_LUT_2C0C 16'h2C0B
`define CUBE_LUT_2C0D 16'h2C0C
`define CUBE_LUT_2C0E 16'h2C0D
`define CUBE_LUT_2C0F 16'h2C0E
`define CUBE_LUT_2C10 16'h2C0F
`define CUBE_LUT_2C11 16'h2C10
`define CUBE_LUT_2C12 16'h2C11
`define CUBE_LUT_2C13 16'h2C12
`define CUBE_LUT_2C14 16'h2C13
`define CUBE_LUT_2C15 16'h2C14
`define CUBE_LUT_2C16 16'h2C15
`define CUBE_LUT_2C17 16'h2C16
`define CUBE_LUT_2C18 16'h2C17
`define CUBE_LUT_2C19 16'h2C18
`define CUBE_LUT_2C1A 16'h2C19
`define CUBE_LUT_2C1B 16'h2C1A
`define CUBE_LUT_2C1C 16'h2C1B
`define CUBE_LUT_2C1D 16'h2C1C
`define CUBE_LUT_2C1E 16'h2C1D
`define CUBE_LUT_2C1F 16'h2C1E
`define CUBE_LUT_2C20 16'h2C1F
`define CUBE_LUT_2C21 16'h2C20
`define CUBE_LUT_2C22 16'h2C21
`define CUBE_LUT_2C23 16'h2C22
`define CUBE_LUT_2C24 16'h2C23
`define CUBE_LUT_2C25 16'h2C24
`define CUBE_LUT_2C26 16'h2C25
`define CUBE_LUT_2C27 16'h2C26
`define CUBE_LUT_2C28 16'h2C27
`define CUBE_LUT_2C29 16'h2C28
`define CUBE_LUT_2C2A 16'h2C28
`define CUBE_LUT_2C2B 16'h2C29
`define CUBE_LUT_2C2C 16'h2C2A
`define CUBE_LUT_2C2D 16'h2C2B
`define CUBE_LUT_2C2E 16'h2C2C
`define CUBE_LUT_2C2F 16'h2C2D
`define CUBE_LUT_2C30 16'h2C2E
`define CUBE_LUT_2C31 16'h2C2F
`define CUBE_LUT_2C32 16'h2C30
`define CUBE_LUT_2C33 16'h2C31
`define CUBE_LUT_2C34 16'h2C32
`define CUBE_LUT_2C35 16'h2C33
`define CUBE_LUT_2C36 16'h2C34
`define CUBE_LUT_2C37 16'h2C35
`define CUBE_LUT_2C38 16'h2C36
`define CUBE_LUT_2C39 16'h2C37
`define CUBE_LUT_2C3A 16'h2C38
`define CUBE_LUT_2C3B 16'h2C39
`define CUBE_LUT_2C3C 16'h2C3A
`define CUBE_LUT_2C3D 16'h2C3B
`define CUBE_LUT_2C3E 16'h2C3C
`define CUBE_LUT_2C3F 16'h2C3D
`define CUBE_LUT_2C40 16'h2C3E
`define CUBE_LUT_2C41 16'h2C3F
`define CUBE_LUT_2C42 16'h2C40
`define CUBE_LUT_2C43 16'h2C41
`define CUBE_LUT_2C44 16'h2C42
`define CUBE_LUT_2C45 16'h2C43
`define CUBE_LUT_2C46 16'h2C44
`define CUBE_LUT_2C47 16'h2C45
`define CUBE_LUT_2C48 16'h2C46
`define CUBE_LUT_2C49 16'h2C47
`define CUBE_LUT_2C4A 16'h2C48
`define CUBE_LUT_2C4B 16'h2C49
`define CUBE_LUT_2C4C 16'h2C4A
`define CUBE_LUT_2C4D 16'h2C4B
`define CUBE_LUT_2C4E 16'h2C4C
`define CUBE_LUT_2C4F 16'h2C4D
`define CUBE_LUT_2C50 16'h2C4E
`define CUBE_LUT_2C51 16'h2C4F
`define CUBE_LUT_2C52 16'h2C50
`define CUBE_LUT_2C53 16'h2C51
`define CUBE_LUT_2C54 16'h2C52
`define CUBE_LUT_2C55 16'h2C53
`define CUBE_LUT_2C56 16'h2C54
`define CUBE_LUT_2C57 16'h2C55
`define CUBE_LUT_2C58 16'h2C56
`define CUBE_LUT_2C59 16'h2C57
`define CUBE_LUT_2C5A 16'h2C58
`define CUBE_LUT_2C5B 16'h2C59
`define CUBE_LUT_2C5C 16'h2C5A
`define CUBE_LUT_2C5D 16'h2C5B
`define CUBE_LUT_2C5E 16'h2C5C
`define CUBE_LUT_2C5F 16'h2C5D
`define CUBE_LUT_2C60 16'h2C5E
`define CUBE_LUT_2C61 16'h2C5F
`define CUBE_LUT_2C62 16'h2C60
`define CUBE_LUT_2C63 16'h2C61
`define CUBE_LUT_2C64 16'h2C62
`define CUBE_LUT_2C65 16'h2C63
`define CUBE_LUT_2C66 16'h2C64
`define CUBE_LUT_2C67 16'h2C65
`define CUBE_LUT_2C68 16'h2C66
`define CUBE_LUT_2C69 16'h2C67
`define CUBE_LUT_2C6A 16'h2C68
`define CUBE_LUT_2C6B 16'h2C69
`define CUBE_LUT_2C6C 16'h2C6A
`define CUBE_LUT_2C6D 16'h2C6B
`define CUBE_LUT_2C6E 16'h2C6C
`define CUBE_LUT_2C6F 16'h2C6D
`define CUBE_LUT_2C70 16'h2C6E
`define CUBE_LUT_2C71 16'h2C6F
`define CUBE_LUT_2C72 16'h2C70
`define CUBE_LUT_2C73 16'h2C71
`define CUBE_LUT_2C74 16'h2C72
`define CUBE_LUT_2C75 16'h2C73
`define CUBE_LUT_2C76 16'h2C74
`define CUBE_LUT_2C77 16'h2C75
`define CUBE_LUT_2C78 16'h2C76
`define CUBE_LUT_2C79 16'h2C77
`define CUBE_LUT_2C7A 16'h2C78
`define CUBE_LUT_2C7B 16'h2C79
`define CUBE_LUT_2C7C 16'h2C7A
`define CUBE_LUT_2C7D 16'h2C7B
`define CUBE_LUT_2C7E 16'h2C7C
`define CUBE_LUT_2C7F 16'h2C7D
`define CUBE_LUT_2C80 16'h2C7E
`define CUBE_LUT_2C81 16'h2C7F
`define CUBE_LUT_2C82 16'h2C80
`define CUBE_LUT_2C83 16'h2C81
`define CUBE_LUT_2C84 16'h2C82
`define CUBE_LUT_2C85 16'h2C83
`define CUBE_LUT_2C86 16'h2C84
`define CUBE_LUT_2C87 16'h2C85
`define CUBE_LUT_2C88 16'h2C86
`define CUBE_LUT_2C89 16'h2C87
`define CUBE_LUT_2C8A 16'h2C88
`define CUBE_LUT_2C8B 16'h2C89
`define CUBE_LUT_2C8C 16'h2C8A
`define CUBE_LUT_2C8D 16'h2C8B
`define CUBE_LUT_2C8E 16'h2C8C
`define CUBE_LUT_2C8F 16'h2C8D
`define CUBE_LUT_2C90 16'h2C8E
`define CUBE_LUT_2C91 16'h2C8F
`define CUBE_LUT_2C92 16'h2C90
`define CUBE_LUT_2C93 16'h2C91
`define CUBE_LUT_2C94 16'h2C92
`define CUBE_LUT_2C95 16'h2C93
`define CUBE_LUT_2C96 16'h2C94
`define CUBE_LUT_2C97 16'h2C95
`define CUBE_LUT_2C98 16'h2C96
`define CUBE_LUT_2C99 16'h2C97
`define CUBE_LUT_2C9A 16'h2C98
`define CUBE_LUT_2C9B 16'h2C99
`define CUBE_LUT_2C9C 16'h2C9A
`define CUBE_LUT_2C9D 16'h2C9B
`define CUBE_LUT_2C9E 16'h2C9C
`define CUBE_LUT_2C9F 16'h2C9D
`define CUBE_LUT_2CA0 16'h2C9E
`define CUBE_LUT_2CA1 16'h2C9F
`define CUBE_LUT_2CA2 16'h2CA0
`define CUBE_LUT_2CA3 16'h2CA1
`define CUBE_LUT_2CA4 16'h2CA2
`define CUBE_LUT_2CA5 16'h2CA3
`define CUBE_LUT_2CA6 16'h2CA4
`define CUBE_LUT_2CA7 16'h2CA5
`define CUBE_LUT_2CA8 16'h2CA6
`define CUBE_LUT_2CA9 16'h2CA7
`define CUBE_LUT_2CAA 16'h2CA8
`define CUBE_LUT_2CAB 16'h2CA9
`define CUBE_LUT_2CAC 16'h2CAA
`define CUBE_LUT_2CAD 16'h2CAB
`define CUBE_LUT_2CAE 16'h2CAC
`define CUBE_LUT_2CAF 16'h2CAD
`define CUBE_LUT_2CB0 16'h2CAE
`define CUBE_LUT_2CB1 16'h2CAF
`define CUBE_LUT_2CB2 16'h2CB0
`define CUBE_LUT_2CB3 16'h2CB1
`define CUBE_LUT_2CB4 16'h2CB2
`define CUBE_LUT_2CB5 16'h2CB3
`define CUBE_LUT_2CB6 16'h2CB4
`define CUBE_LUT_2CB7 16'h2CB5
`define CUBE_LUT_2CB8 16'h2CB6
`define CUBE_LUT_2CB9 16'h2CB7
`define CUBE_LUT_2CBA 16'h2CB8
`define CUBE_LUT_2CBB 16'h2CB9
`define CUBE_LUT_2CBC 16'h2CBA
`define CUBE_LUT_2CBD 16'h2CBB
`define CUBE_LUT_2CBE 16'h2CBC
`define CUBE_LUT_2CBF 16'h2CBD
`define CUBE_LUT_2CC0 16'h2CBE
`define CUBE_LUT_2CC1 16'h2CBF
`define CUBE_LUT_2CC2 16'h2CC0
`define CUBE_LUT_2CC3 16'h2CC1
`define CUBE_LUT_2CC4 16'h2CC2
`define CUBE_LUT_2CC5 16'h2CC3
`define CUBE_LUT_2CC6 16'h2CC4
`define CUBE_LUT_2CC7 16'h2CC5
`define CUBE_LUT_2CC8 16'h2CC6
`define CUBE_LUT_2CC9 16'h2CC7
`define CUBE_LUT_2CCA 16'h2CC8
`define CUBE_LUT_2CCB 16'h2CC9
`define CUBE_LUT_2CCC 16'h2CCA
`define CUBE_LUT_2CCD 16'h2CCB
`define CUBE_LUT_2CCE 16'h2CCC
`define CUBE_LUT_2CCF 16'h2CCD
`define CUBE_LUT_2CD0 16'h2CCE
`define CUBE_LUT_2CD1 16'h2CCF
`define CUBE_LUT_2CD2 16'h2CD0
`define CUBE_LUT_2CD3 16'h2CD1
`define CUBE_LUT_2CD4 16'h2CD2
`define CUBE_LUT_2CD5 16'h2CD3
`define CUBE_LUT_2CD6 16'h2CD4
`define CUBE_LUT_2CD7 16'h2CD5
`define CUBE_LUT_2CD8 16'h2CD6
`define CUBE_LUT_2CD9 16'h2CD7
`define CUBE_LUT_2CDA 16'h2CD8
`define CUBE_LUT_2CDB 16'h2CD9
`define CUBE_LUT_2CDC 16'h2CDA
`define CUBE_LUT_2CDD 16'h2CDB
`define CUBE_LUT_2CDE 16'h2CDC
`define CUBE_LUT_2CDF 16'h2CDD
`define CUBE_LUT_2CE0 16'h2CDE
`define CUBE_LUT_2CE1 16'h2CDF
`define CUBE_LUT_2CE2 16'h2CE0
`define CUBE_LUT_2CE3 16'h2CE1
`define CUBE_LUT_2CE4 16'h2CE2
`define CUBE_LUT_2CE5 16'h2CE3
`define CUBE_LUT_2CE6 16'h2CE4
`define CUBE_LUT_2CE7 16'h2CE5
`define CUBE_LUT_2CE8 16'h2CE6
`define CUBE_LUT_2CE9 16'h2CE7
`define CUBE_LUT_2CEA 16'h2CE8
`define CUBE_LUT_2CEB 16'h2CE9
`define CUBE_LUT_2CEC 16'h2CEA
`define CUBE_LUT_2CED 16'h2CEB
`define CUBE_LUT_2CEE 16'h2CEC
`define CUBE_LUT_2CEF 16'h2CED
`define CUBE_LUT_2CF0 16'h2CED
`define CUBE_LUT_2CF1 16'h2CEE
`define CUBE_LUT_2CF2 16'h2CEF
`define CUBE_LUT_2CF3 16'h2CF0
`define CUBE_LUT_2CF4 16'h2CF1
`define CUBE_LUT_2CF5 16'h2CF2
`define CUBE_LUT_2CF6 16'h2CF3
`define CUBE_LUT_2CF7 16'h2CF4
`define CUBE_LUT_2CF8 16'h2CF5
`define CUBE_LUT_2CF9 16'h2CF6
`define CUBE_LUT_2CFA 16'h2CF7
`define CUBE_LUT_2CFB 16'h2CF8
`define CUBE_LUT_2CFC 16'h2CF9
`define CUBE_LUT_2CFD 16'h2CFA
`define CUBE_LUT_2CFE 16'h2CFB
`define CUBE_LUT_2CFF 16'h2CFC
`define CUBE_LUT_2D00 16'h2CFD
`define CUBE_LUT_2D01 16'h2CFE
`define CUBE_LUT_2D02 16'h2CFF
`define CUBE_LUT_2D03 16'h2D00
`define CUBE_LUT_2D04 16'h2D01
`define CUBE_LUT_2D05 16'h2D02
`define CUBE_LUT_2D06 16'h2D03
`define CUBE_LUT_2D07 16'h2D04
`define CUBE_LUT_2D08 16'h2D05
`define CUBE_LUT_2D09 16'h2D06
`define CUBE_LUT_2D0A 16'h2D07
`define CUBE_LUT_2D0B 16'h2D08
`define CUBE_LUT_2D0C 16'h2D09
`define CUBE_LUT_2D0D 16'h2D0A
`define CUBE_LUT_2D0E 16'h2D0B
`define CUBE_LUT_2D0F 16'h2D0C
`define CUBE_LUT_2D10 16'h2D0D
`define CUBE_LUT_2D11 16'h2D0E
`define CUBE_LUT_2D12 16'h2D0F
`define CUBE_LUT_2D13 16'h2D10
`define CUBE_LUT_2D14 16'h2D11
`define CUBE_LUT_2D15 16'h2D12
`define CUBE_LUT_2D16 16'h2D13
`define CUBE_LUT_2D17 16'h2D14
`define CUBE_LUT_2D18 16'h2D15
`define CUBE_LUT_2D19 16'h2D16
`define CUBE_LUT_2D1A 16'h2D17
`define CUBE_LUT_2D1B 16'h2D18
`define CUBE_LUT_2D1C 16'h2D19
`define CUBE_LUT_2D1D 16'h2D1A
`define CUBE_LUT_2D1E 16'h2D1B
`define CUBE_LUT_2D1F 16'h2D1C
`define CUBE_LUT_2D20 16'h2D1D
`define CUBE_LUT_2D21 16'h2D1E
`define CUBE_LUT_2D22 16'h2D1F
`define CUBE_LUT_2D23 16'h2D20
`define CUBE_LUT_2D24 16'h2D21
`define CUBE_LUT_2D25 16'h2D22
`define CUBE_LUT_2D26 16'h2D23
`define CUBE_LUT_2D27 16'h2D24
`define CUBE_LUT_2D28 16'h2D25
`define CUBE_LUT_2D29 16'h2D26
`define CUBE_LUT_2D2A 16'h2D27
`define CUBE_LUT_2D2B 16'h2D28
`define CUBE_LUT_2D2C 16'h2D29
`define CUBE_LUT_2D2D 16'h2D2A
`define CUBE_LUT_2D2E 16'h2D2B
`define CUBE_LUT_2D2F 16'h2D2C
`define CUBE_LUT_2D30 16'h2D2D
`define CUBE_LUT_2D31 16'h2D2E
`define CUBE_LUT_2D32 16'h2D2F
`define CUBE_LUT_2D33 16'h2D30
`define CUBE_LUT_2D34 16'h2D31
`define CUBE_LUT_2D35 16'h2D32
`define CUBE_LUT_2D36 16'h2D33
`define CUBE_LUT_2D37 16'h2D34
`define CUBE_LUT_2D38 16'h2D35
`define CUBE_LUT_2D39 16'h2D36
`define CUBE_LUT_2D3A 16'h2D37
`define CUBE_LUT_2D3B 16'h2D38
`define CUBE_LUT_2D3C 16'h2D39
`define CUBE_LUT_2D3D 16'h2D3A
`define CUBE_LUT_2D3E 16'h2D3B
`define CUBE_LUT_2D3F 16'h2D3C
`define CUBE_LUT_2D40 16'h2D3D
`define CUBE_LUT_2D41 16'h2D3E
`define CUBE_LUT_2D42 16'h2D3F
`define CUBE_LUT_2D43 16'h2D40
`define CUBE_LUT_2D44 16'h2D41
`define CUBE_LUT_2D45 16'h2D42
`define CUBE_LUT_2D46 16'h2D43
`define CUBE_LUT_2D47 16'h2D44
`define CUBE_LUT_2D48 16'h2D45
`define CUBE_LUT_2D49 16'h2D46
`define CUBE_LUT_2D4A 16'h2D47
`define CUBE_LUT_2D4B 16'h2D48
`define CUBE_LUT_2D4C 16'h2D49
`define CUBE_LUT_2D4D 16'h2D4A
`define CUBE_LUT_2D4E 16'h2D4B
`define CUBE_LUT_2D4F 16'h2D4C
`define CUBE_LUT_2D50 16'h2D4D
`define CUBE_LUT_2D51 16'h2D4E
`define CUBE_LUT_2D52 16'h2D4F
`define CUBE_LUT_2D53 16'h2D50
`define CUBE_LUT_2D54 16'h2D51
`define CUBE_LUT_2D55 16'h2D52
`define CUBE_LUT_2D56 16'h2D53
`define CUBE_LUT_2D57 16'h2D54
`define CUBE_LUT_2D58 16'h2D55
`define CUBE_LUT_2D59 16'h2D56
`define CUBE_LUT_2D5A 16'h2D57
`define CUBE_LUT_2D5B 16'h2D58
`define CUBE_LUT_2D5C 16'h2D59
`define CUBE_LUT_2D5D 16'h2D5A
`define CUBE_LUT_2D5E 16'h2D5B
`define CUBE_LUT_2D5F 16'h2D5C
`define CUBE_LUT_2D60 16'h2D5D
`define CUBE_LUT_2D61 16'h2D5E
`define CUBE_LUT_2D62 16'h2D5F
`define CUBE_LUT_2D63 16'h2D60
`define CUBE_LUT_2D64 16'h2D61
`define CUBE_LUT_2D65 16'h2D62
`define CUBE_LUT_2D66 16'h2D63
`define CUBE_LUT_2D67 16'h2D64
`define CUBE_LUT_2D68 16'h2D65
`define CUBE_LUT_2D69 16'h2D66
`define CUBE_LUT_2D6A 16'h2D67
`define CUBE_LUT_2D6B 16'h2D68
`define CUBE_LUT_2D6C 16'h2D69
`define CUBE_LUT_2D6D 16'h2D6A
`define CUBE_LUT_2D6E 16'h2D6B
`define CUBE_LUT_2D6F 16'h2D6C
`define CUBE_LUT_2D70 16'h2D6D
`define CUBE_LUT_2D71 16'h2D6E
`define CUBE_LUT_2D72 16'h2D6F
`define CUBE_LUT_2D73 16'h2D70
`define CUBE_LUT_2D74 16'h2D71
`define CUBE_LUT_2D75 16'h2D72
`define CUBE_LUT_2D76 16'h2D73
`define CUBE_LUT_2D77 16'h2D74
`define CUBE_LUT_2D78 16'h2D75
`define CUBE_LUT_2D79 16'h2D76
`define CUBE_LUT_2D7A 16'h2D77
`define CUBE_LUT_2D7B 16'h2D78
`define CUBE_LUT_2D7C 16'h2D79
`define CUBE_LUT_2D7D 16'h2D7A
`define CUBE_LUT_2D7E 16'h2D7B
`define CUBE_LUT_2D7F 16'h2D7C
`define CUBE_LUT_2D80 16'h2D7D
`define CUBE_LUT_2D81 16'h2D7E
`define CUBE_LUT_2D82 16'h2D7F
`define CUBE_LUT_2D83 16'h2D80
`define CUBE_LUT_2D84 16'h2D81
`define CUBE_LUT_2D85 16'h2D82
`define CUBE_LUT_2D86 16'h2D82
`define CUBE_LUT_2D87 16'h2D83
`define CUBE_LUT_2D88 16'h2D84
`define CUBE_LUT_2D89 16'h2D85
`define CUBE_LUT_2D8A 16'h2D86
`define CUBE_LUT_2D8B 16'h2D87
`define CUBE_LUT_2D8C 16'h2D88
`define CUBE_LUT_2D8D 16'h2D89
`define CUBE_LUT_2D8E 16'h2D8A
`define CUBE_LUT_2D8F 16'h2D8B
`define CUBE_LUT_2D90 16'h2D8C
`define CUBE_LUT_2D91 16'h2D8D
`define CUBE_LUT_2D92 16'h2D8E
`define CUBE_LUT_2D93 16'h2D8F
`define CUBE_LUT_2D94 16'h2D90
`define CUBE_LUT_2D95 16'h2D91
`define CUBE_LUT_2D96 16'h2D92
`define CUBE_LUT_2D97 16'h2D93
`define CUBE_LUT_2D98 16'h2D94
`define CUBE_LUT_2D99 16'h2D95
`define CUBE_LUT_2D9A 16'h2D96
`define CUBE_LUT_2D9B 16'h2D97
`define CUBE_LUT_2D9C 16'h2D98
`define CUBE_LUT_2D9D 16'h2D99
`define CUBE_LUT_2D9E 16'h2D9A
`define CUBE_LUT_2D9F 16'h2D9B
`define CUBE_LUT_2DA0 16'h2D9C
`define CUBE_LUT_2DA1 16'h2D9D
`define CUBE_LUT_2DA2 16'h2D9E
`define CUBE_LUT_2DA3 16'h2D9F
`define CUBE_LUT_2DA4 16'h2DA0
`define CUBE_LUT_2DA5 16'h2DA1
`define CUBE_LUT_2DA6 16'h2DA2
`define CUBE_LUT_2DA7 16'h2DA3
`define CUBE_LUT_2DA8 16'h2DA4
`define CUBE_LUT_2DA9 16'h2DA5
`define CUBE_LUT_2DAA 16'h2DA6
`define CUBE_LUT_2DAB 16'h2DA7
`define CUBE_LUT_2DAC 16'h2DA8
`define CUBE_LUT_2DAD 16'h2DA9
`define CUBE_LUT_2DAE 16'h2DAA
`define CUBE_LUT_2DAF 16'h2DAB
`define CUBE_LUT_2DB0 16'h2DAC
`define CUBE_LUT_2DB1 16'h2DAD
`define CUBE_LUT_2DB2 16'h2DAE
`define CUBE_LUT_2DB3 16'h2DAF
`define CUBE_LUT_2DB4 16'h2DB0
`define CUBE_LUT_2DB5 16'h2DB1
`define CUBE_LUT_2DB6 16'h2DB2
`define CUBE_LUT_2DB7 16'h2DB3
`define CUBE_LUT_2DB8 16'h2DB4
`define CUBE_LUT_2DB9 16'h2DB5
`define CUBE_LUT_2DBA 16'h2DB6
`define CUBE_LUT_2DBB 16'h2DB7
`define CUBE_LUT_2DBC 16'h2DB8
`define CUBE_LUT_2DBD 16'h2DB9
`define CUBE_LUT_2DBE 16'h2DBA
`define CUBE_LUT_2DBF 16'h2DBB
`define CUBE_LUT_2DC0 16'h2DBC
`define CUBE_LUT_2DC1 16'h2DBD
`define CUBE_LUT_2DC2 16'h2DBE
`define CUBE_LUT_2DC3 16'h2DBF
`define CUBE_LUT_2DC4 16'h2DC0
`define CUBE_LUT_2DC5 16'h2DC1
`define CUBE_LUT_2DC6 16'h2DC2
`define CUBE_LUT_2DC7 16'h2DC3
`define CUBE_LUT_2DC8 16'h2DC4
`define CUBE_LUT_2DC9 16'h2DC5
`define CUBE_LUT_2DCA 16'h2DC6
`define CUBE_LUT_2DCB 16'h2DC7
`define CUBE_LUT_2DCC 16'h2DC8
`define CUBE_LUT_2DCD 16'h2DC9
`define CUBE_LUT_2DCE 16'h2DCA
`define CUBE_LUT_2DCF 16'h2DCB
`define CUBE_LUT_2DD0 16'h2DCC
`define CUBE_LUT_2DD1 16'h2DCD
`define CUBE_LUT_2DD2 16'h2DCE
`define CUBE_LUT_2DD3 16'h2DCF
`define CUBE_LUT_2DD4 16'h2DD0
`define CUBE_LUT_2DD5 16'h2DD1
`define CUBE_LUT_2DD6 16'h2DD2
`define CUBE_LUT_2DD7 16'h2DD3
`define CUBE_LUT_2DD8 16'h2DD4
`define CUBE_LUT_2DD9 16'h2DD5
`define CUBE_LUT_2DDA 16'h2DD6
`define CUBE_LUT_2DDB 16'h2DD7
`define CUBE_LUT_2DDC 16'h2DD8
`define CUBE_LUT_2DDD 16'h2DD9
`define CUBE_LUT_2DDE 16'h2DDA
`define CUBE_LUT_2DDF 16'h2DDB
`define CUBE_LUT_2DE0 16'h2DDC
`define CUBE_LUT_2DE1 16'h2DDD
`define CUBE_LUT_2DE2 16'h2DDE
`define CUBE_LUT_2DE3 16'h2DDF
`define CUBE_LUT_2DE4 16'h2DE0
`define CUBE_LUT_2DE5 16'h2DE1
`define CUBE_LUT_2DE6 16'h2DE2
`define CUBE_LUT_2DE7 16'h2DE3
`define CUBE_LUT_2DE8 16'h2DE4
`define CUBE_LUT_2DE9 16'h2DE5
`define CUBE_LUT_2DEA 16'h2DE6
`define CUBE_LUT_2DEB 16'h2DE7
`define CUBE_LUT_2DEC 16'h2DE8
`define CUBE_LUT_2DED 16'h2DE9
`define CUBE_LUT_2DEE 16'h2DEA
`define CUBE_LUT_2DEF 16'h2DEB
`define CUBE_LUT_2DF0 16'h2DEC
`define CUBE_LUT_2DF1 16'h2DED
`define CUBE_LUT_2DF2 16'h2DEE
`define CUBE_LUT_2DF3 16'h2DEF
`define CUBE_LUT_2DF4 16'h2DF0
`define CUBE_LUT_2DF5 16'h2DF1
`define CUBE_LUT_2DF6 16'h2DF2
`define CUBE_LUT_2DF7 16'h2DF3
`define CUBE_LUT_2DF8 16'h2DF4
`define CUBE_LUT_2DF9 16'h2DF5
`define CUBE_LUT_2DFA 16'h2DF6
`define CUBE_LUT_2DFB 16'h2DF7
`define CUBE_LUT_2DFC 16'h2DF8
`define CUBE_LUT_2DFD 16'h2DF9
`define CUBE_LUT_2DFE 16'h2DFA
`define CUBE_LUT_2DFF 16'h2DFB
`define CUBE_LUT_2E00 16'h2DFC
`define CUBE_LUT_2E01 16'h2DFD
`define CUBE_LUT_2E02 16'h2DFD
`define CUBE_LUT_2E03 16'h2DFE
`define CUBE_LUT_2E04 16'h2DFF
`define CUBE_LUT_2E05 16'h2E00
`define CUBE_LUT_2E06 16'h2E01
`define CUBE_LUT_2E07 16'h2E02
`define CUBE_LUT_2E08 16'h2E03
`define CUBE_LUT_2E09 16'h2E04
`define CUBE_LUT_2E0A 16'h2E05
`define CUBE_LUT_2E0B 16'h2E06
`define CUBE_LUT_2E0C 16'h2E07
`define CUBE_LUT_2E0D 16'h2E08
`define CUBE_LUT_2E0E 16'h2E09
`define CUBE_LUT_2E0F 16'h2E0A
`define CUBE_LUT_2E10 16'h2E0B
`define CUBE_LUT_2E11 16'h2E0C
`define CUBE_LUT_2E12 16'h2E0D
`define CUBE_LUT_2E13 16'h2E0E
`define CUBE_LUT_2E14 16'h2E0F
`define CUBE_LUT_2E15 16'h2E10
`define CUBE_LUT_2E16 16'h2E11
`define CUBE_LUT_2E17 16'h2E12
`define CUBE_LUT_2E18 16'h2E13
`define CUBE_LUT_2E19 16'h2E14
`define CUBE_LUT_2E1A 16'h2E15
`define CUBE_LUT_2E1B 16'h2E16
`define CUBE_LUT_2E1C 16'h2E17
`define CUBE_LUT_2E1D 16'h2E18
`define CUBE_LUT_2E1E 16'h2E19
`define CUBE_LUT_2E1F 16'h2E1A
`define CUBE_LUT_2E20 16'h2E1B
`define CUBE_LUT_2E21 16'h2E1C
`define CUBE_LUT_2E22 16'h2E1D
`define CUBE_LUT_2E23 16'h2E1E
`define CUBE_LUT_2E24 16'h2E1F
`define CUBE_LUT_2E25 16'h2E20
`define CUBE_LUT_2E26 16'h2E21
`define CUBE_LUT_2E27 16'h2E22
`define CUBE_LUT_2E28 16'h2E23
`define CUBE_LUT_2E29 16'h2E24
`define CUBE_LUT_2E2A 16'h2E25
`define CUBE_LUT_2E2B 16'h2E26
`define CUBE_LUT_2E2C 16'h2E27
`define CUBE_LUT_2E2D 16'h2E28
`define CUBE_LUT_2E2E 16'h2E29
`define CUBE_LUT_2E2F 16'h2E2A
`define CUBE_LUT_2E30 16'h2E2B
`define CUBE_LUT_2E31 16'h2E2C
`define CUBE_LUT_2E32 16'h2E2D
`define CUBE_LUT_2E33 16'h2E2E
`define CUBE_LUT_2E34 16'h2E2F
`define CUBE_LUT_2E35 16'h2E30
`define CUBE_LUT_2E36 16'h2E31
`define CUBE_LUT_2E37 16'h2E32
`define CUBE_LUT_2E38 16'h2E33
`define CUBE_LUT_2E39 16'h2E34
`define CUBE_LUT_2E3A 16'h2E35
`define CUBE_LUT_2E3B 16'h2E36
`define CUBE_LUT_2E3C 16'h2E37
`define CUBE_LUT_2E3D 16'h2E38
`define CUBE_LUT_2E3E 16'h2E39
`define CUBE_LUT_2E3F 16'h2E3A
`define CUBE_LUT_2E40 16'h2E3B
`define CUBE_LUT_2E41 16'h2E3C
`define CUBE_LUT_2E42 16'h2E3D
`define CUBE_LUT_2E43 16'h2E3E
`define CUBE_LUT_2E44 16'h2E3F
`define CUBE_LUT_2E45 16'h2E40
`define CUBE_LUT_2E46 16'h2E41
`define CUBE_LUT_2E47 16'h2E42
`define CUBE_LUT_2E48 16'h2E43
`define CUBE_LUT_2E49 16'h2E44
`define CUBE_LUT_2E4A 16'h2E45
`define CUBE_LUT_2E4B 16'h2E46
`define CUBE_LUT_2E4C 16'h2E47
`define CUBE_LUT_2E4D 16'h2E48
`define CUBE_LUT_2E4E 16'h2E49
`define CUBE_LUT_2E4F 16'h2E4A
`define CUBE_LUT_2E50 16'h2E4B
`define CUBE_LUT_2E51 16'h2E4C
`define CUBE_LUT_2E52 16'h2E4D
`define CUBE_LUT_2E53 16'h2E4E
`define CUBE_LUT_2E54 16'h2E4F
`define CUBE_LUT_2E55 16'h2E50
`define CUBE_LUT_2E56 16'h2E51
`define CUBE_LUT_2E57 16'h2E52
`define CUBE_LUT_2E58 16'h2E53
`define CUBE_LUT_2E59 16'h2E54
`define CUBE_LUT_2E5A 16'h2E55
`define CUBE_LUT_2E5B 16'h2E56
`define CUBE_LUT_2E5C 16'h2E57
`define CUBE_LUT_2E5D 16'h2E58
`define CUBE_LUT_2E5E 16'h2E59
`define CUBE_LUT_2E5F 16'h2E5A
`define CUBE_LUT_2E60 16'h2E5B
`define CUBE_LUT_2E61 16'h2E5C
`define CUBE_LUT_2E62 16'h2E5D
`define CUBE_LUT_2E63 16'h2E5E
`define CUBE_LUT_2E64 16'h2E5F
`define CUBE_LUT_2E65 16'h2E60
`define CUBE_LUT_2E66 16'h2E61
`define CUBE_LUT_2E67 16'h2E62
`define CUBE_LUT_2E68 16'h2E63
`define CUBE_LUT_2E69 16'h2E64
`define CUBE_LUT_2E6A 16'h2E65
`define CUBE_LUT_2E6B 16'h2E66
`define CUBE_LUT_2E6C 16'h2E67
`define CUBE_LUT_2E6D 16'h2E67
`define CUBE_LUT_2E6E 16'h2E68
`define CUBE_LUT_2E6F 16'h2E69
`define CUBE_LUT_2E70 16'h2E6A
`define CUBE_LUT_2E71 16'h2E6B
`define CUBE_LUT_2E72 16'h2E6C
`define CUBE_LUT_2E73 16'h2E6D
`define CUBE_LUT_2E74 16'h2E6E
`define CUBE_LUT_2E75 16'h2E6F
`define CUBE_LUT_2E76 16'h2E70
`define CUBE_LUT_2E77 16'h2E71
`define CUBE_LUT_2E78 16'h2E72
`define CUBE_LUT_2E79 16'h2E73
`define CUBE_LUT_2E7A 16'h2E74
`define CUBE_LUT_2E7B 16'h2E75
`define CUBE_LUT_2E7C 16'h2E76
`define CUBE_LUT_2E7D 16'h2E77
`define CUBE_LUT_2E7E 16'h2E78
`define CUBE_LUT_2E7F 16'h2E79
`define CUBE_LUT_2E80 16'h2E7A
`define CUBE_LUT_2E81 16'h2E7B
`define CUBE_LUT_2E82 16'h2E7C
`define CUBE_LUT_2E83 16'h2E7D
`define CUBE_LUT_2E84 16'h2E7E
`define CUBE_LUT_2E85 16'h2E7F
`define CUBE_LUT_2E86 16'h2E80
`define CUBE_LUT_2E87 16'h2E81
`define CUBE_LUT_2E88 16'h2E82
`define CUBE_LUT_2E89 16'h2E83
`define CUBE_LUT_2E8A 16'h2E84
`define CUBE_LUT_2E8B 16'h2E85
`define CUBE_LUT_2E8C 16'h2E86
`define CUBE_LUT_2E8D 16'h2E87
`define CUBE_LUT_2E8E 16'h2E88
`define CUBE_LUT_2E8F 16'h2E89
`define CUBE_LUT_2E90 16'h2E8A
`define CUBE_LUT_2E91 16'h2E8B
`define CUBE_LUT_2E92 16'h2E8C
`define CUBE_LUT_2E93 16'h2E8D
`define CUBE_LUT_2E94 16'h2E8E
`define CUBE_LUT_2E95 16'h2E8F
`define CUBE_LUT_2E96 16'h2E90
`define CUBE_LUT_2E97 16'h2E91
`define CUBE_LUT_2E98 16'h2E92
`define CUBE_LUT_2E99 16'h2E93
`define CUBE_LUT_2E9A 16'h2E94
`define CUBE_LUT_2E9B 16'h2E95
`define CUBE_LUT_2E9C 16'h2E96
`define CUBE_LUT_2E9D 16'h2E97
`define CUBE_LUT_2E9E 16'h2E98
`define CUBE_LUT_2E9F 16'h2E99
`define CUBE_LUT_2EA0 16'h2E9A
`define CUBE_LUT_2EA1 16'h2E9B
`define CUBE_LUT_2EA2 16'h2E9C
`define CUBE_LUT_2EA3 16'h2E9D
`define CUBE_LUT_2EA4 16'h2E9E
`define CUBE_LUT_2EA5 16'h2E9F
`define CUBE_LUT_2EA6 16'h2EA0
`define CUBE_LUT_2EA7 16'h2EA1
`define CUBE_LUT_2EA8 16'h2EA2
`define CUBE_LUT_2EA9 16'h2EA3
`define CUBE_LUT_2EAA 16'h2EA4
`define CUBE_LUT_2EAB 16'h2EA5
`define CUBE_LUT_2EAC 16'h2EA6
`define CUBE_LUT_2EAD 16'h2EA7
`define CUBE_LUT_2EAE 16'h2EA8
`define CUBE_LUT_2EAF 16'h2EA9
`define CUBE_LUT_2EB0 16'h2EAA
`define CUBE_LUT_2EB1 16'h2EAB
`define CUBE_LUT_2EB2 16'h2EAC
`define CUBE_LUT_2EB3 16'h2EAD
`define CUBE_LUT_2EB4 16'h2EAE
`define CUBE_LUT_2EB5 16'h2EAF
`define CUBE_LUT_2EB6 16'h2EB0
`define CUBE_LUT_2EB7 16'h2EB1
`define CUBE_LUT_2EB8 16'h2EB2
`define CUBE_LUT_2EB9 16'h2EB3
`define CUBE_LUT_2EBA 16'h2EB4
`define CUBE_LUT_2EBB 16'h2EB5
`define CUBE_LUT_2EBC 16'h2EB6
`define CUBE_LUT_2EBD 16'h2EB7
`define CUBE_LUT_2EBE 16'h2EB8
`define CUBE_LUT_2EBF 16'h2EB9
`define CUBE_LUT_2EC0 16'h2EBA
`define CUBE_LUT_2EC1 16'h2EBB
`define CUBE_LUT_2EC2 16'h2EBC
`define CUBE_LUT_2EC3 16'h2EBD
`define CUBE_LUT_2EC4 16'h2EBE
`define CUBE_LUT_2EC5 16'h2EBF
`define CUBE_LUT_2EC6 16'h2EC0
`define CUBE_LUT_2EC7 16'h2EC1
`define CUBE_LUT_2EC8 16'h2EC2
`define CUBE_LUT_2EC9 16'h2EC3
`define CUBE_LUT_2ECA 16'h2EC4
`define CUBE_LUT_2ECB 16'h2EC4
`define CUBE_LUT_2ECC 16'h2EC5
`define CUBE_LUT_2ECD 16'h2EC6
`define CUBE_LUT_2ECE 16'h2EC7
`define CUBE_LUT_2ECF 16'h2EC8
`define CUBE_LUT_2ED0 16'h2EC9
`define CUBE_LUT_2ED1 16'h2ECA
`define CUBE_LUT_2ED2 16'h2ECB
`define CUBE_LUT_2ED3 16'h2ECC
`define CUBE_LUT_2ED4 16'h2ECD
`define CUBE_LUT_2ED5 16'h2ECE
`define CUBE_LUT_2ED6 16'h2ECF
`define CUBE_LUT_2ED7 16'h2ED0
`define CUBE_LUT_2ED8 16'h2ED1
`define CUBE_LUT_2ED9 16'h2ED2
`define CUBE_LUT_2EDA 16'h2ED3
`define CUBE_LUT_2EDB 16'h2ED4
`define CUBE_LUT_2EDC 16'h2ED5
`define CUBE_LUT_2EDD 16'h2ED6
`define CUBE_LUT_2EDE 16'h2ED7
`define CUBE_LUT_2EDF 16'h2ED8
`define CUBE_LUT_2EE0 16'h2ED9
`define CUBE_LUT_2EE1 16'h2EDA
`define CUBE_LUT_2EE2 16'h2EDB
`define CUBE_LUT_2EE3 16'h2EDC
`define CUBE_LUT_2EE4 16'h2EDD
`define CUBE_LUT_2EE5 16'h2EDE
`define CUBE_LUT_2EE6 16'h2EDF
`define CUBE_LUT_2EE7 16'h2EE0
`define CUBE_LUT_2EE8 16'h2EE1
`define CUBE_LUT_2EE9 16'h2EE2
`define CUBE_LUT_2EEA 16'h2EE3
`define CUBE_LUT_2EEB 16'h2EE4
`define CUBE_LUT_2EEC 16'h2EE5
`define CUBE_LUT_2EED 16'h2EE6
`define CUBE_LUT_2EEE 16'h2EE7
`define CUBE_LUT_2EEF 16'h2EE8
`define CUBE_LUT_2EF0 16'h2EE9
`define CUBE_LUT_2EF1 16'h2EEA
`define CUBE_LUT_2EF2 16'h2EEB
`define CUBE_LUT_2EF3 16'h2EEC
`define CUBE_LUT_2EF4 16'h2EED
`define CUBE_LUT_2EF5 16'h2EEE
`define CUBE_LUT_2EF6 16'h2EEF
`define CUBE_LUT_2EF7 16'h2EF0
`define CUBE_LUT_2EF8 16'h2EF1
`define CUBE_LUT_2EF9 16'h2EF2
`define CUBE_LUT_2EFA 16'h2EF3
`define CUBE_LUT_2EFB 16'h2EF4
`define CUBE_LUT_2EFC 16'h2EF5
`define CUBE_LUT_2EFD 16'h2EF6
`define CUBE_LUT_2EFE 16'h2EF7
`define CUBE_LUT_2EFF 16'h2EF8
`define CUBE_LUT_2F00 16'h2EF9
`define CUBE_LUT_2F01 16'h2EFA
`define CUBE_LUT_2F02 16'h2EFB
`define CUBE_LUT_2F03 16'h2EFC
`define CUBE_LUT_2F04 16'h2EFD
`define CUBE_LUT_2F05 16'h2EFE
`define CUBE_LUT_2F06 16'h2EFF
`define CUBE_LUT_2F07 16'h2F00
`define CUBE_LUT_2F08 16'h2F01
`define CUBE_LUT_2F09 16'h2F02
`define CUBE_LUT_2F0A 16'h2F03
`define CUBE_LUT_2F0B 16'h2F04
`define CUBE_LUT_2F0C 16'h2F05
`define CUBE_LUT_2F0D 16'h2F06
`define CUBE_LUT_2F0E 16'h2F07
`define CUBE_LUT_2F0F 16'h2F08
`define CUBE_LUT_2F10 16'h2F09
`define CUBE_LUT_2F11 16'h2F0A
`define CUBE_LUT_2F12 16'h2F0B
`define CUBE_LUT_2F13 16'h2F0C
`define CUBE_LUT_2F14 16'h2F0D
`define CUBE_LUT_2F15 16'h2F0E
`define CUBE_LUT_2F16 16'h2F0F
`define CUBE_LUT_2F17 16'h2F10
`define CUBE_LUT_2F18 16'h2F11
`define CUBE_LUT_2F19 16'h2F12
`define CUBE_LUT_2F1A 16'h2F13
`define CUBE_LUT_2F1B 16'h2F14
`define CUBE_LUT_2F1C 16'h2F15
`define CUBE_LUT_2F1D 16'h2F16
`define CUBE_LUT_2F1E 16'h2F17
`define CUBE_LUT_2F1F 16'h2F18
`define CUBE_LUT_2F20 16'h2F19
`define CUBE_LUT_2F21 16'h2F19
`define CUBE_LUT_2F22 16'h2F1A
`define CUBE_LUT_2F23 16'h2F1B
`define CUBE_LUT_2F24 16'h2F1C
`define CUBE_LUT_2F25 16'h2F1D
`define CUBE_LUT_2F26 16'h2F1E
`define CUBE_LUT_2F27 16'h2F1F
`define CUBE_LUT_2F28 16'h2F20
`define CUBE_LUT_2F29 16'h2F21
`define CUBE_LUT_2F2A 16'h2F22
`define CUBE_LUT_2F2B 16'h2F23
`define CUBE_LUT_2F2C 16'h2F24
`define CUBE_LUT_2F2D 16'h2F25
`define CUBE_LUT_2F2E 16'h2F26
`define CUBE_LUT_2F2F 16'h2F27
`define CUBE_LUT_2F30 16'h2F28
`define CUBE_LUT_2F31 16'h2F29
`define CUBE_LUT_2F32 16'h2F2A
`define CUBE_LUT_2F33 16'h2F2B
`define CUBE_LUT_2F34 16'h2F2C
`define CUBE_LUT_2F35 16'h2F2D
`define CUBE_LUT_2F36 16'h2F2E
`define CUBE_LUT_2F37 16'h2F2F
`define CUBE_LUT_2F38 16'h2F30
`define CUBE_LUT_2F39 16'h2F31
`define CUBE_LUT_2F3A 16'h2F32
`define CUBE_LUT_2F3B 16'h2F33
`define CUBE_LUT_2F3C 16'h2F34
`define CUBE_LUT_2F3D 16'h2F35
`define CUBE_LUT_2F3E 16'h2F36
`define CUBE_LUT_2F3F 16'h2F37
`define CUBE_LUT_2F40 16'h2F38
`define CUBE_LUT_2F41 16'h2F39
`define CUBE_LUT_2F42 16'h2F3A
`define CUBE_LUT_2F43 16'h2F3B
`define CUBE_LUT_2F44 16'h2F3C
`define CUBE_LUT_2F45 16'h2F3D
`define CUBE_LUT_2F46 16'h2F3E
`define CUBE_LUT_2F47 16'h2F3F
`define CUBE_LUT_2F48 16'h2F40
`define CUBE_LUT_2F49 16'h2F41
`define CUBE_LUT_2F4A 16'h2F42
`define CUBE_LUT_2F4B 16'h2F43
`define CUBE_LUT_2F4C 16'h2F44
`define CUBE_LUT_2F4D 16'h2F45
`define CUBE_LUT_2F4E 16'h2F46
`define CUBE_LUT_2F4F 16'h2F47
`define CUBE_LUT_2F50 16'h2F48
`define CUBE_LUT_2F51 16'h2F49
`define CUBE_LUT_2F52 16'h2F4A
`define CUBE_LUT_2F53 16'h2F4B
`define CUBE_LUT_2F54 16'h2F4C
`define CUBE_LUT_2F55 16'h2F4D
`define CUBE_LUT_2F56 16'h2F4E
`define CUBE_LUT_2F57 16'h2F4F
`define CUBE_LUT_2F58 16'h2F50
`define CUBE_LUT_2F59 16'h2F51
`define CUBE_LUT_2F5A 16'h2F52
`define CUBE_LUT_2F5B 16'h2F53
`define CUBE_LUT_2F5C 16'h2F54
`define CUBE_LUT_2F5D 16'h2F55
`define CUBE_LUT_2F5E 16'h2F56
`define CUBE_LUT_2F5F 16'h2F57
`define CUBE_LUT_2F60 16'h2F58
`define CUBE_LUT_2F61 16'h2F59
`define CUBE_LUT_2F62 16'h2F5A
`define CUBE_LUT_2F63 16'h2F5B
`define CUBE_LUT_2F64 16'h2F5C
`define CUBE_LUT_2F65 16'h2F5D
`define CUBE_LUT_2F66 16'h2F5E
`define CUBE_LUT_2F67 16'h2F5F
`define CUBE_LUT_2F68 16'h2F60
`define CUBE_LUT_2F69 16'h2F61
`define CUBE_LUT_2F6A 16'h2F62
`define CUBE_LUT_2F6B 16'h2F63
`define CUBE_LUT_2F6C 16'h2F64
`define CUBE_LUT_2F6D 16'h2F65
`define CUBE_LUT_2F6E 16'h2F66
`define CUBE_LUT_2F6F 16'h2F66
`define CUBE_LUT_2F70 16'h2F67
`define CUBE_LUT_2F71 16'h2F68
`define CUBE_LUT_2F72 16'h2F69
`define CUBE_LUT_2F73 16'h2F6A
`define CUBE_LUT_2F74 16'h2F6B
`define CUBE_LUT_2F75 16'h2F6C
`define CUBE_LUT_2F76 16'h2F6D
`define CUBE_LUT_2F77 16'h2F6E
`define CUBE_LUT_2F78 16'h2F6F
`define CUBE_LUT_2F79 16'h2F70
`define CUBE_LUT_2F7A 16'h2F71
`define CUBE_LUT_2F7B 16'h2F72
`define CUBE_LUT_2F7C 16'h2F73
`define CUBE_LUT_2F7D 16'h2F74
`define CUBE_LUT_2F7E 16'h2F75
`define CUBE_LUT_2F7F 16'h2F76
`define CUBE_LUT_2F80 16'h2F77
`define CUBE_LUT_2F81 16'h2F78
`define CUBE_LUT_2F82 16'h2F79
`define CUBE_LUT_2F83 16'h2F7A
`define CUBE_LUT_2F84 16'h2F7B
`define CUBE_LUT_2F85 16'h2F7C
`define CUBE_LUT_2F86 16'h2F7D
`define CUBE_LUT_2F87 16'h2F7E
`define CUBE_LUT_2F88 16'h2F7F
`define CUBE_LUT_2F89 16'h2F80
`define CUBE_LUT_2F8A 16'h2F81
`define CUBE_LUT_2F8B 16'h2F82
`define CUBE_LUT_2F8C 16'h2F83
`define CUBE_LUT_2F8D 16'h2F84
`define CUBE_LUT_2F8E 16'h2F85
`define CUBE_LUT_2F8F 16'h2F86
`define CUBE_LUT_2F90 16'h2F87
`define CUBE_LUT_2F91 16'h2F88
`define CUBE_LUT_2F92 16'h2F89
`define CUBE_LUT_2F93 16'h2F8A
`define CUBE_LUT_2F94 16'h2F8B
`define CUBE_LUT_2F95 16'h2F8C
`define CUBE_LUT_2F96 16'h2F8D
`define CUBE_LUT_2F97 16'h2F8E
`define CUBE_LUT_2F98 16'h2F8F
`define CUBE_LUT_2F99 16'h2F90
`define CUBE_LUT_2F9A 16'h2F91
`define CUBE_LUT_2F9B 16'h2F92
`define CUBE_LUT_2F9C 16'h2F93
`define CUBE_LUT_2F9D 16'h2F94
`define CUBE_LUT_2F9E 16'h2F95
`define CUBE_LUT_2F9F 16'h2F96
`define CUBE_LUT_2FA0 16'h2F97
`define CUBE_LUT_2FA1 16'h2F98
`define CUBE_LUT_2FA2 16'h2F99
`define CUBE_LUT_2FA3 16'h2F9A
`define CUBE_LUT_2FA4 16'h2F9B
`define CUBE_LUT_2FA5 16'h2F9C
`define CUBE_LUT_2FA6 16'h2F9D
`define CUBE_LUT_2FA7 16'h2F9E
`define CUBE_LUT_2FA8 16'h2F9F
`define CUBE_LUT_2FA9 16'h2FA0
`define CUBE_LUT_2FAA 16'h2FA1
`define CUBE_LUT_2FAB 16'h2FA2
`define CUBE_LUT_2FAC 16'h2FA3
`define CUBE_LUT_2FAD 16'h2FA4
`define CUBE_LUT_2FAE 16'h2FA5
`define CUBE_LUT_2FAF 16'h2FA6
`define CUBE_LUT_2FB0 16'h2FA7
`define CUBE_LUT_2FB1 16'h2FA8
`define CUBE_LUT_2FB2 16'h2FA9
`define CUBE_LUT_2FB3 16'h2FAA
`define CUBE_LUT_2FB4 16'h2FAB
`define CUBE_LUT_2FB5 16'h2FAC
`define CUBE_LUT_2FB6 16'h2FAD
`define CUBE_LUT_2FB7 16'h2FAD
`define CUBE_LUT_2FB8 16'h2FAE
`define CUBE_LUT_2FB9 16'h2FAF
`define CUBE_LUT_2FBA 16'h2FB0
`define CUBE_LUT_2FBB 16'h2FB1
`define CUBE_LUT_2FBC 16'h2FB2
`define CUBE_LUT_2FBD 16'h2FB3
`define CUBE_LUT_2FBE 16'h2FB4
`define CUBE_LUT_2FBF 16'h2FB5
`define CUBE_LUT_2FC0 16'h2FB6
`define CUBE_LUT_2FC1 16'h2FB7
`define CUBE_LUT_2FC2 16'h2FB8
`define CUBE_LUT_2FC3 16'h2FB9
`define CUBE_LUT_2FC4 16'h2FBA
`define CUBE_LUT_2FC5 16'h2FBB
`define CUBE_LUT_2FC6 16'h2FBC
`define CUBE_LUT_2FC7 16'h2FBD
`define CUBE_LUT_2FC8 16'h2FBE
`define CUBE_LUT_2FC9 16'h2FBF
`define CUBE_LUT_2FCA 16'h2FC0
`define CUBE_LUT_2FCB 16'h2FC1
`define CUBE_LUT_2FCC 16'h2FC2
`define CUBE_LUT_2FCD 16'h2FC3
`define CUBE_LUT_2FCE 16'h2FC4
`define CUBE_LUT_2FCF 16'h2FC5
`define CUBE_LUT_2FD0 16'h2FC6
`define CUBE_LUT_2FD1 16'h2FC7
`define CUBE_LUT_2FD2 16'h2FC8
`define CUBE_LUT_2FD3 16'h2FC9
`define CUBE_LUT_2FD4 16'h2FCA
`define CUBE_LUT_2FD5 16'h2FCB
`define CUBE_LUT_2FD6 16'h2FCC
`define CUBE_LUT_2FD7 16'h2FCD
`define CUBE_LUT_2FD8 16'h2FCE
`define CUBE_LUT_2FD9 16'h2FCF
`define CUBE_LUT_2FDA 16'h2FD0
`define CUBE_LUT_2FDB 16'h2FD1
`define CUBE_LUT_2FDC 16'h2FD2
`define CUBE_LUT_2FDD 16'h2FD3
`define CUBE_LUT_2FDE 16'h2FD4
`define CUBE_LUT_2FDF 16'h2FD5
`define CUBE_LUT_2FE0 16'h2FD6
`define CUBE_LUT_2FE1 16'h2FD7
`define CUBE_LUT_2FE2 16'h2FD8
`define CUBE_LUT_2FE3 16'h2FD9
`define CUBE_LUT_2FE4 16'h2FDA
`define CUBE_LUT_2FE5 16'h2FDB
`define CUBE_LUT_2FE6 16'h2FDC
`define CUBE_LUT_2FE7 16'h2FDD
`define CUBE_LUT_2FE8 16'h2FDE
`define CUBE_LUT_2FE9 16'h2FDF
`define CUBE_LUT_2FEA 16'h2FE0
`define CUBE_LUT_2FEB 16'h2FE1
`define CUBE_LUT_2FEC 16'h2FE2
`define CUBE_LUT_2FED 16'h2FE3
`define CUBE_LUT_2FEE 16'h2FE4
`define CUBE_LUT_2FEF 16'h2FE5
`define CUBE_LUT_2FF0 16'h2FE6
`define CUBE_LUT_2FF1 16'h2FE7
`define CUBE_LUT_2FF2 16'h2FE8
`define CUBE_LUT_2FF3 16'h2FE9
`define CUBE_LUT_2FF4 16'h2FEA
`define CUBE_LUT_2FF5 16'h2FEB
`define CUBE_LUT_2FF6 16'h2FEC
`define CUBE_LUT_2FF7 16'h2FED
`define CUBE_LUT_2FF8 16'h2FEE
`define CUBE_LUT_2FF9 16'h2FEF
`define CUBE_LUT_2FFA 16'h2FEF
`define CUBE_LUT_2FFB 16'h2FF0
`define CUBE_LUT_2FFC 16'h2FF1
`define CUBE_LUT_2FFD 16'h2FF2
`define CUBE_LUT_2FFE 16'h2FF3
`define CUBE_LUT_2FFF 16'h2FF4
`define CUBE_LUT_3000 16'h2FF5
`define CUBE_LUT_3001 16'h2FF7
`define CUBE_LUT_3002 16'h2FF9
`define CUBE_LUT_3003 16'h2FFB
`define CUBE_LUT_3004 16'h2FFD
`define CUBE_LUT_3005 16'h2FFF
`define CUBE_LUT_3006 16'h3001
`define CUBE_LUT_3007 16'h3002
`define CUBE_LUT_3008 16'h3003
`define CUBE_LUT_3009 16'h3004
`define CUBE_LUT_300A 16'h3005
`define CUBE_LUT_300B 16'h3006
`define CUBE_LUT_300C 16'h3007
`define CUBE_LUT_300D 16'h3007
`define CUBE_LUT_300E 16'h3008
`define CUBE_LUT_300F 16'h3009
`define CUBE_LUT_3010 16'h300A
`define CUBE_LUT_3011 16'h300B
`define CUBE_LUT_3012 16'h300C
`define CUBE_LUT_3013 16'h300D
`define CUBE_LUT_3014 16'h300E
`define CUBE_LUT_3015 16'h300F
`define CUBE_LUT_3016 16'h3010
`define CUBE_LUT_3017 16'h3011
`define CUBE_LUT_3018 16'h3012
`define CUBE_LUT_3019 16'h3013
`define CUBE_LUT_301A 16'h3014
`define CUBE_LUT_301B 16'h3015
`define CUBE_LUT_301C 16'h3016
`define CUBE_LUT_301D 16'h3017
`define CUBE_LUT_301E 16'h3018
`define CUBE_LUT_301F 16'h3019
`define CUBE_LUT_3020 16'h301A
`define CUBE_LUT_3021 16'h301B
`define CUBE_LUT_3022 16'h301C
`define CUBE_LUT_3023 16'h301D
`define CUBE_LUT_3024 16'h301E
`define CUBE_LUT_3025 16'h301F
`define CUBE_LUT_3026 16'h3020
`define CUBE_LUT_3027 16'h3021
`define CUBE_LUT_3028 16'h3022
`define CUBE_LUT_3029 16'h3023
`define CUBE_LUT_302A 16'h3024
`define CUBE_LUT_302B 16'h3025
`define CUBE_LUT_302C 16'h3026
`define CUBE_LUT_302D 16'h3027
`define CUBE_LUT_302E 16'h3028
`define CUBE_LUT_302F 16'h3029
`define CUBE_LUT_3030 16'h302A
`define CUBE_LUT_3031 16'h302B
`define CUBE_LUT_3032 16'h302C
`define CUBE_LUT_3033 16'h302D
`define CUBE_LUT_3034 16'h302E
`define CUBE_LUT_3035 16'h302F
`define CUBE_LUT_3036 16'h3030
`define CUBE_LUT_3037 16'h3031
`define CUBE_LUT_3038 16'h3032
`define CUBE_LUT_3039 16'h3033
`define CUBE_LUT_303A 16'h3034
`define CUBE_LUT_303B 16'h3035
`define CUBE_LUT_303C 16'h3036
`define CUBE_LUT_303D 16'h3037
`define CUBE_LUT_303E 16'h3038
`define CUBE_LUT_303F 16'h3039
`define CUBE_LUT_3040 16'h303A
`define CUBE_LUT_3041 16'h303B
`define CUBE_LUT_3042 16'h303C
`define CUBE_LUT_3043 16'h303D
`define CUBE_LUT_3044 16'h303E
`define CUBE_LUT_3045 16'h303F
`define CUBE_LUT_3046 16'h3040
`define CUBE_LUT_3047 16'h3041
`define CUBE_LUT_3048 16'h3042
`define CUBE_LUT_3049 16'h3042
`define CUBE_LUT_304A 16'h3043
`define CUBE_LUT_304B 16'h3044
`define CUBE_LUT_304C 16'h3045
`define CUBE_LUT_304D 16'h3046
`define CUBE_LUT_304E 16'h3047
`define CUBE_LUT_304F 16'h3048
`define CUBE_LUT_3050 16'h3049
`define CUBE_LUT_3051 16'h304A
`define CUBE_LUT_3052 16'h304B
`define CUBE_LUT_3053 16'h304C
`define CUBE_LUT_3054 16'h304D
`define CUBE_LUT_3055 16'h304E
`define CUBE_LUT_3056 16'h304F
`define CUBE_LUT_3057 16'h3050
`define CUBE_LUT_3058 16'h3051
`define CUBE_LUT_3059 16'h3052
`define CUBE_LUT_305A 16'h3053
`define CUBE_LUT_305B 16'h3054
`define CUBE_LUT_305C 16'h3055
`define CUBE_LUT_305D 16'h3056
`define CUBE_LUT_305E 16'h3057
`define CUBE_LUT_305F 16'h3058
`define CUBE_LUT_3060 16'h3059
`define CUBE_LUT_3061 16'h305A
`define CUBE_LUT_3062 16'h305B
`define CUBE_LUT_3063 16'h305C
`define CUBE_LUT_3064 16'h305D
`define CUBE_LUT_3065 16'h305E
`define CUBE_LUT_3066 16'h305F
`define CUBE_LUT_3067 16'h3060
`define CUBE_LUT_3068 16'h3061
`define CUBE_LUT_3069 16'h3062
`define CUBE_LUT_306A 16'h3063
`define CUBE_LUT_306B 16'h3064
`define CUBE_LUT_306C 16'h3065
`define CUBE_LUT_306D 16'h3066
`define CUBE_LUT_306E 16'h3067
`define CUBE_LUT_306F 16'h3068
`define CUBE_LUT_3070 16'h3069
`define CUBE_LUT_3071 16'h306A
`define CUBE_LUT_3072 16'h306B
`define CUBE_LUT_3073 16'h306C
`define CUBE_LUT_3074 16'h306D
`define CUBE_LUT_3075 16'h306E
`define CUBE_LUT_3076 16'h306F
`define CUBE_LUT_3077 16'h3070
`define CUBE_LUT_3078 16'h3071
`define CUBE_LUT_3079 16'h3072
`define CUBE_LUT_307A 16'h3073
`define CUBE_LUT_307B 16'h3074
`define CUBE_LUT_307C 16'h3075
`define CUBE_LUT_307D 16'h3076
`define CUBE_LUT_307E 16'h3077
`define CUBE_LUT_307F 16'h3077
`define CUBE_LUT_3080 16'h3078
`define CUBE_LUT_3081 16'h3079
`define CUBE_LUT_3082 16'h307A
`define CUBE_LUT_3083 16'h307B
`define CUBE_LUT_3084 16'h307C
`define CUBE_LUT_3085 16'h307D
`define CUBE_LUT_3086 16'h307E
`define CUBE_LUT_3087 16'h307F
`define CUBE_LUT_3088 16'h3080
`define CUBE_LUT_3089 16'h3081
`define CUBE_LUT_308A 16'h3082
`define CUBE_LUT_308B 16'h3083
`define CUBE_LUT_308C 16'h3084
`define CUBE_LUT_308D 16'h3085
`define CUBE_LUT_308E 16'h3086
`define CUBE_LUT_308F 16'h3087
`define CUBE_LUT_3090 16'h3088
`define CUBE_LUT_3091 16'h3089
`define CUBE_LUT_3092 16'h308A
`define CUBE_LUT_3093 16'h308B
`define CUBE_LUT_3094 16'h308C
`define CUBE_LUT_3095 16'h308D
`define CUBE_LUT_3096 16'h308E
`define CUBE_LUT_3097 16'h308F
`define CUBE_LUT_3098 16'h3090
`define CUBE_LUT_3099 16'h3091
`define CUBE_LUT_309A 16'h3092
`define CUBE_LUT_309B 16'h3093
`define CUBE_LUT_309C 16'h3094
`define CUBE_LUT_309D 16'h3095
`define CUBE_LUT_309E 16'h3096
`define CUBE_LUT_309F 16'h3097
`define CUBE_LUT_30A0 16'h3098
`define CUBE_LUT_30A1 16'h3099
`define CUBE_LUT_30A2 16'h309A
`define CUBE_LUT_30A3 16'h309B
`define CUBE_LUT_30A4 16'h309C
`define CUBE_LUT_30A5 16'h309D
`define CUBE_LUT_30A6 16'h309E
`define CUBE_LUT_30A7 16'h309F
`define CUBE_LUT_30A8 16'h30A0
`define CUBE_LUT_30A9 16'h30A1
`define CUBE_LUT_30AA 16'h30A2
`define CUBE_LUT_30AB 16'h30A3
`define CUBE_LUT_30AC 16'h30A4
`define CUBE_LUT_30AD 16'h30A5
`define CUBE_LUT_30AE 16'h30A6
`define CUBE_LUT_30AF 16'h30A7
`define CUBE_LUT_30B0 16'h30A7
`define CUBE_LUT_30B1 16'h30A8
`define CUBE_LUT_30B2 16'h30A9
`define CUBE_LUT_30B3 16'h30AA
`define CUBE_LUT_30B4 16'h30AB
`define CUBE_LUT_30B5 16'h30AC
`define CUBE_LUT_30B6 16'h30AD
`define CUBE_LUT_30B7 16'h30AE
`define CUBE_LUT_30B8 16'h30AF
`define CUBE_LUT_30B9 16'h30B0
`define CUBE_LUT_30BA 16'h30B1
`define CUBE_LUT_30BB 16'h30B2
`define CUBE_LUT_30BC 16'h30B3
`define CUBE_LUT_30BD 16'h30B4
`define CUBE_LUT_30BE 16'h30B5
`define CUBE_LUT_30BF 16'h30B6
`define CUBE_LUT_30C0 16'h30B7
`define CUBE_LUT_30C1 16'h30B8
`define CUBE_LUT_30C2 16'h30B9
`define CUBE_LUT_30C3 16'h30BA
`define CUBE_LUT_30C4 16'h30BB
`define CUBE_LUT_30C5 16'h30BC
`define CUBE_LUT_30C6 16'h30BD
`define CUBE_LUT_30C7 16'h30BE
`define CUBE_LUT_30C8 16'h30BF
`define CUBE_LUT_30C9 16'h30C0
`define CUBE_LUT_30CA 16'h30C1
`define CUBE_LUT_30CB 16'h30C2
`define CUBE_LUT_30CC 16'h30C3
`define CUBE_LUT_30CD 16'h30C4
`define CUBE_LUT_30CE 16'h30C5
`define CUBE_LUT_30CF 16'h30C6
`define CUBE_LUT_30D0 16'h30C7
`define CUBE_LUT_30D1 16'h30C8
`define CUBE_LUT_30D2 16'h30C9
`define CUBE_LUT_30D3 16'h30CA
`define CUBE_LUT_30D4 16'h30CB
`define CUBE_LUT_30D5 16'h30CC
`define CUBE_LUT_30D6 16'h30CD
`define CUBE_LUT_30D7 16'h30CE
`define CUBE_LUT_30D8 16'h30CF
`define CUBE_LUT_30D9 16'h30D0
`define CUBE_LUT_30DA 16'h30D1
`define CUBE_LUT_30DB 16'h30D2
`define CUBE_LUT_30DC 16'h30D3
`define CUBE_LUT_30DD 16'h30D4
`define CUBE_LUT_30DE 16'h30D4
`define CUBE_LUT_30DF 16'h30D5
`define CUBE_LUT_30E0 16'h30D6
`define CUBE_LUT_30E1 16'h30D7
`define CUBE_LUT_30E2 16'h30D8
`define CUBE_LUT_30E3 16'h30D9
`define CUBE_LUT_30E4 16'h30DA
`define CUBE_LUT_30E5 16'h30DB
`define CUBE_LUT_30E6 16'h30DC
`define CUBE_LUT_30E7 16'h30DD
`define CUBE_LUT_30E8 16'h30DE
`define CUBE_LUT_30E9 16'h30DF
`define CUBE_LUT_30EA 16'h30E0
`define CUBE_LUT_30EB 16'h30E1
`define CUBE_LUT_30EC 16'h30E2
`define CUBE_LUT_30ED 16'h30E3
`define CUBE_LUT_30EE 16'h30E4
`define CUBE_LUT_30EF 16'h30E5
`define CUBE_LUT_30F0 16'h30E6
`define CUBE_LUT_30F1 16'h30E7
`define CUBE_LUT_30F2 16'h30E8
`define CUBE_LUT_30F3 16'h30E9
`define CUBE_LUT_30F4 16'h30EA
`define CUBE_LUT_30F5 16'h30EB
`define CUBE_LUT_30F6 16'h30EC
`define CUBE_LUT_30F7 16'h30ED
`define CUBE_LUT_30F8 16'h30EE
`define CUBE_LUT_30F9 16'h30EF
`define CUBE_LUT_30FA 16'h30F0
`define CUBE_LUT_30FB 16'h30F1
`define CUBE_LUT_30FC 16'h30F2
`define CUBE_LUT_30FD 16'h30F3
`define CUBE_LUT_30FE 16'h30F4
`define CUBE_LUT_30FF 16'h30F5
`define CUBE_LUT_3100 16'h30F6
`define CUBE_LUT_3101 16'h30F7
`define CUBE_LUT_3102 16'h30F8
`define CUBE_LUT_3103 16'h30F9
`define CUBE_LUT_3104 16'h30FA
`define CUBE_LUT_3105 16'h30FB
`define CUBE_LUT_3106 16'h30FC
`define CUBE_LUT_3107 16'h30FD
`define CUBE_LUT_3108 16'h30FD
`define CUBE_LUT_3109 16'h30FE
`define CUBE_LUT_310A 16'h30FF
`define CUBE_LUT_310B 16'h3100
`define CUBE_LUT_310C 16'h3101
`define CUBE_LUT_310D 16'h3102
`define CUBE_LUT_310E 16'h3103
`define CUBE_LUT_310F 16'h3104
`define CUBE_LUT_3110 16'h3105
`define CUBE_LUT_3111 16'h3106
`define CUBE_LUT_3112 16'h3107
`define CUBE_LUT_3113 16'h3108
`define CUBE_LUT_3114 16'h3109
`define CUBE_LUT_3115 16'h310A
`define CUBE_LUT_3116 16'h310B
`define CUBE_LUT_3117 16'h310C
`define CUBE_LUT_3118 16'h310D
`define CUBE_LUT_3119 16'h310E
`define CUBE_LUT_311A 16'h310F
`define CUBE_LUT_311B 16'h3110
`define CUBE_LUT_311C 16'h3111
`define CUBE_LUT_311D 16'h3112
`define CUBE_LUT_311E 16'h3113
`define CUBE_LUT_311F 16'h3114
`define CUBE_LUT_3120 16'h3115
`define CUBE_LUT_3121 16'h3116
`define CUBE_LUT_3122 16'h3117
`define CUBE_LUT_3123 16'h3118
`define CUBE_LUT_3124 16'h3119
`define CUBE_LUT_3125 16'h311A
`define CUBE_LUT_3126 16'h311B
`define CUBE_LUT_3127 16'h311C
`define CUBE_LUT_3128 16'h311D
`define CUBE_LUT_3129 16'h311E
`define CUBE_LUT_312A 16'h311F
`define CUBE_LUT_312B 16'h3120
`define CUBE_LUT_312C 16'h3121
`define CUBE_LUT_312D 16'h3122
`define CUBE_LUT_312E 16'h3123
`define CUBE_LUT_312F 16'h3124
`define CUBE_LUT_3130 16'h3124
`define CUBE_LUT_3131 16'h3125
`define CUBE_LUT_3132 16'h3126
`define CUBE_LUT_3133 16'h3127
`define CUBE_LUT_3134 16'h3128
`define CUBE_LUT_3135 16'h3129
`define CUBE_LUT_3136 16'h312A
`define CUBE_LUT_3137 16'h312B
`define CUBE_LUT_3138 16'h312C
`define CUBE_LUT_3139 16'h312D
`define CUBE_LUT_313A 16'h312E
`define CUBE_LUT_313B 16'h312F
`define CUBE_LUT_313C 16'h3130
`define CUBE_LUT_313D 16'h3131
`define CUBE_LUT_313E 16'h3132
`define CUBE_LUT_313F 16'h3133
`define CUBE_LUT_3140 16'h3134
`define CUBE_LUT_3141 16'h3135
`define CUBE_LUT_3142 16'h3136
`define CUBE_LUT_3143 16'h3137
`define CUBE_LUT_3144 16'h3138
`define CUBE_LUT_3145 16'h3139
`define CUBE_LUT_3146 16'h313A
`define CUBE_LUT_3147 16'h313B
`define CUBE_LUT_3148 16'h313C
`define CUBE_LUT_3149 16'h313D
`define CUBE_LUT_314A 16'h313E
`define CUBE_LUT_314B 16'h313F
`define CUBE_LUT_314C 16'h3140
`define CUBE_LUT_314D 16'h3141
`define CUBE_LUT_314E 16'h3142
`define CUBE_LUT_314F 16'h3143
`define CUBE_LUT_3150 16'h3144
`define CUBE_LUT_3151 16'h3145
`define CUBE_LUT_3152 16'h3146
`define CUBE_LUT_3153 16'h3147
`define CUBE_LUT_3154 16'h3148
`define CUBE_LUT_3155 16'h3149
`define CUBE_LUT_3156 16'h3149
`define CUBE_LUT_3157 16'h314A
`define CUBE_LUT_3158 16'h314B
`define CUBE_LUT_3159 16'h314C
`define CUBE_LUT_315A 16'h314D
`define CUBE_LUT_315B 16'h314E
`define CUBE_LUT_315C 16'h314F
`define CUBE_LUT_315D 16'h3150
`define CUBE_LUT_315E 16'h3151
`define CUBE_LUT_315F 16'h3152
`define CUBE_LUT_3160 16'h3153
`define CUBE_LUT_3161 16'h3154
`define CUBE_LUT_3162 16'h3155
`define CUBE_LUT_3163 16'h3156
`define CUBE_LUT_3164 16'h3157
`define CUBE_LUT_3165 16'h3158
`define CUBE_LUT_3166 16'h3159
`define CUBE_LUT_3167 16'h315A
`define CUBE_LUT_3168 16'h315B
`define CUBE_LUT_3169 16'h315C
`define CUBE_LUT_316A 16'h315D
`define CUBE_LUT_316B 16'h315E
`define CUBE_LUT_316C 16'h315F
`define CUBE_LUT_316D 16'h3160
`define CUBE_LUT_316E 16'h3161
`define CUBE_LUT_316F 16'h3162
`define CUBE_LUT_3170 16'h3163
`define CUBE_LUT_3171 16'h3164
`define CUBE_LUT_3172 16'h3165
`define CUBE_LUT_3173 16'h3166
`define CUBE_LUT_3174 16'h3167
`define CUBE_LUT_3175 16'h3168
`define CUBE_LUT_3176 16'h3169
`define CUBE_LUT_3177 16'h316A
`define CUBE_LUT_3178 16'h316B
`define CUBE_LUT_3179 16'h316B
`define CUBE_LUT_317A 16'h316C
`define CUBE_LUT_317B 16'h316D
`define CUBE_LUT_317C 16'h316E
`define CUBE_LUT_317D 16'h316F
`define CUBE_LUT_317E 16'h3170
`define CUBE_LUT_317F 16'h3171
`define CUBE_LUT_3180 16'h3172
`define CUBE_LUT_3181 16'h3173
`define CUBE_LUT_3182 16'h3174
`define CUBE_LUT_3183 16'h3175
`define CUBE_LUT_3184 16'h3176
`define CUBE_LUT_3185 16'h3177
`define CUBE_LUT_3186 16'h3178
`define CUBE_LUT_3187 16'h3179
`define CUBE_LUT_3188 16'h317A
`define CUBE_LUT_3189 16'h317B
`define CUBE_LUT_318A 16'h317C
`define CUBE_LUT_318B 16'h317D
`define CUBE_LUT_318C 16'h317E
`define CUBE_LUT_318D 16'h317F
`define CUBE_LUT_318E 16'h3180
`define CUBE_LUT_318F 16'h3181
`define CUBE_LUT_3190 16'h3182
`define CUBE_LUT_3191 16'h3183
`define CUBE_LUT_3192 16'h3184
`define CUBE_LUT_3193 16'h3185
`define CUBE_LUT_3194 16'h3186
`define CUBE_LUT_3195 16'h3187
`define CUBE_LUT_3196 16'h3188
`define CUBE_LUT_3197 16'h3189
`define CUBE_LUT_3198 16'h318A
`define CUBE_LUT_3199 16'h318B
`define CUBE_LUT_319A 16'h318C
`define CUBE_LUT_319B 16'h318D
`define CUBE_LUT_319C 16'h318D
`define CUBE_LUT_319D 16'h318E
`define CUBE_LUT_319E 16'h318F
`define CUBE_LUT_319F 16'h3190
`define CUBE_LUT_31A0 16'h3191
`define CUBE_LUT_31A1 16'h3192
`define CUBE_LUT_31A2 16'h3193
`define CUBE_LUT_31A3 16'h3194
`define CUBE_LUT_31A4 16'h3195
`define CUBE_LUT_31A5 16'h3196
`define CUBE_LUT_31A6 16'h3197
`define CUBE_LUT_31A7 16'h3198
`define CUBE_LUT_31A8 16'h3199
`define CUBE_LUT_31A9 16'h319A
`define CUBE_LUT_31AA 16'h319B
`define CUBE_LUT_31AB 16'h319C
`define CUBE_LUT_31AC 16'h319D
`define CUBE_LUT_31AD 16'h319E
`define CUBE_LUT_31AE 16'h319F
`define CUBE_LUT_31AF 16'h31A0
`define CUBE_LUT_31B0 16'h31A1
`define CUBE_LUT_31B1 16'h31A2
`define CUBE_LUT_31B2 16'h31A3
`define CUBE_LUT_31B3 16'h31A4
`define CUBE_LUT_31B4 16'h31A5
`define CUBE_LUT_31B5 16'h31A6
`define CUBE_LUT_31B6 16'h31A7
`define CUBE_LUT_31B7 16'h31A8
`define CUBE_LUT_31B8 16'h31A9
`define CUBE_LUT_31B9 16'h31AA
`define CUBE_LUT_31BA 16'h31AB
`define CUBE_LUT_31BB 16'h31AC
`define CUBE_LUT_31BC 16'h31AC
`define CUBE_LUT_31BD 16'h31AD
`define CUBE_LUT_31BE 16'h31AE
`define CUBE_LUT_31BF 16'h31AF
`define CUBE_LUT_31C0 16'h31B0
`define CUBE_LUT_31C1 16'h31B1
`define CUBE_LUT_31C2 16'h31B2
`define CUBE_LUT_31C3 16'h31B3
`define CUBE_LUT_31C4 16'h31B4
`define CUBE_LUT_31C5 16'h31B5
`define CUBE_LUT_31C6 16'h31B6
`define CUBE_LUT_31C7 16'h31B7
`define CUBE_LUT_31C8 16'h31B8
`define CUBE_LUT_31C9 16'h31B9
`define CUBE_LUT_31CA 16'h31BA
`define CUBE_LUT_31CB 16'h31BB
`define CUBE_LUT_31CC 16'h31BC
`define CUBE_LUT_31CD 16'h31BD
`define CUBE_LUT_31CE 16'h31BE
`define CUBE_LUT_31CF 16'h31BF
`define CUBE_LUT_31D0 16'h31C0
`define CUBE_LUT_31D1 16'h31C1
`define CUBE_LUT_31D2 16'h31C2
`define CUBE_LUT_31D3 16'h31C3
`define CUBE_LUT_31D4 16'h31C4
`define CUBE_LUT_31D5 16'h31C5
`define CUBE_LUT_31D6 16'h31C6
`define CUBE_LUT_31D7 16'h31C7
`define CUBE_LUT_31D8 16'h31C8
`define CUBE_LUT_31D9 16'h31C9
`define CUBE_LUT_31DA 16'h31CA
`define CUBE_LUT_31DB 16'h31CA
`define CUBE_LUT_31DC 16'h31CB
`define CUBE_LUT_31DD 16'h31CC
`define CUBE_LUT_31DE 16'h31CD
`define CUBE_LUT_31DF 16'h31CE
`define CUBE_LUT_31E0 16'h31CF
`define CUBE_LUT_31E1 16'h31D0
`define CUBE_LUT_31E2 16'h31D1
`define CUBE_LUT_31E3 16'h31D2
`define CUBE_LUT_31E4 16'h31D3
`define CUBE_LUT_31E5 16'h31D4
`define CUBE_LUT_31E6 16'h31D5
`define CUBE_LUT_31E7 16'h31D6
`define CUBE_LUT_31E8 16'h31D7
`define CUBE_LUT_31E9 16'h31D8
`define CUBE_LUT_31EA 16'h31D9
`define CUBE_LUT_31EB 16'h31DA
`define CUBE_LUT_31EC 16'h31DB
`define CUBE_LUT_31ED 16'h31DC
`define CUBE_LUT_31EE 16'h31DD
`define CUBE_LUT_31EF 16'h31DE
`define CUBE_LUT_31F0 16'h31DF
`define CUBE_LUT_31F1 16'h31E0
`define CUBE_LUT_31F2 16'h31E1
`define CUBE_LUT_31F3 16'h31E2
`define CUBE_LUT_31F4 16'h31E3
`define CUBE_LUT_31F5 16'h31E4
`define CUBE_LUT_31F6 16'h31E5
`define CUBE_LUT_31F7 16'h31E6
`define CUBE_LUT_31F8 16'h31E7
`define CUBE_LUT_31F9 16'h31E7
`define CUBE_LUT_31FA 16'h31E8
`define CUBE_LUT_31FB 16'h31E9
`define CUBE_LUT_31FC 16'h31EA
`define CUBE_LUT_31FD 16'h31EB
`define CUBE_LUT_31FE 16'h31EC
`define CUBE_LUT_31FF 16'h31ED
`define CUBE_LUT_3200 16'h31EE
`define CUBE_LUT_3201 16'h31EF
`define CUBE_LUT_3202 16'h31F0
`define CUBE_LUT_3203 16'h31F1
`define CUBE_LUT_3204 16'h31F2
`define CUBE_LUT_3205 16'h31F3
`define CUBE_LUT_3206 16'h31F4
`define CUBE_LUT_3207 16'h31F5
`define CUBE_LUT_3208 16'h31F6
`define CUBE_LUT_3209 16'h31F7
`define CUBE_LUT_320A 16'h31F8
`define CUBE_LUT_320B 16'h31F9
`define CUBE_LUT_320C 16'h31FA
`define CUBE_LUT_320D 16'h31FB
`define CUBE_LUT_320E 16'h31FC
`define CUBE_LUT_320F 16'h31FD
`define CUBE_LUT_3210 16'h31FE
`define CUBE_LUT_3211 16'h31FF
`define CUBE_LUT_3212 16'h3200
`define CUBE_LUT_3213 16'h3201
`define CUBE_LUT_3214 16'h3202
`define CUBE_LUT_3215 16'h3203
`define CUBE_LUT_3216 16'h3203
`define CUBE_LUT_3217 16'h3204
`define CUBE_LUT_3218 16'h3205
`define CUBE_LUT_3219 16'h3206
`define CUBE_LUT_321A 16'h3207
`define CUBE_LUT_321B 16'h3208
`define CUBE_LUT_321C 16'h3209
`define CUBE_LUT_321D 16'h320A
`define CUBE_LUT_321E 16'h320B
`define CUBE_LUT_321F 16'h320C
`define CUBE_LUT_3220 16'h320D
`define CUBE_LUT_3221 16'h320E
`define CUBE_LUT_3222 16'h320F
`define CUBE_LUT_3223 16'h3210
`define CUBE_LUT_3224 16'h3211
`define CUBE_LUT_3225 16'h3212
`define CUBE_LUT_3226 16'h3213
`define CUBE_LUT_3227 16'h3214
`define CUBE_LUT_3228 16'h3215
`define CUBE_LUT_3229 16'h3216
`define CUBE_LUT_322A 16'h3217
`define CUBE_LUT_322B 16'h3218
`define CUBE_LUT_322C 16'h3219
`define CUBE_LUT_322D 16'h321A
`define CUBE_LUT_322E 16'h321B
`define CUBE_LUT_322F 16'h321C
`define CUBE_LUT_3230 16'h321D
`define CUBE_LUT_3231 16'h321E
`define CUBE_LUT_3232 16'h321E
`define CUBE_LUT_3233 16'h321F
`define CUBE_LUT_3234 16'h3220
`define CUBE_LUT_3235 16'h3221
`define CUBE_LUT_3236 16'h3222
`define CUBE_LUT_3237 16'h3223
`define CUBE_LUT_3238 16'h3224
`define CUBE_LUT_3239 16'h3225
`define CUBE_LUT_323A 16'h3226
`define CUBE_LUT_323B 16'h3227
`define CUBE_LUT_323C 16'h3228
`define CUBE_LUT_323D 16'h3229
`define CUBE_LUT_323E 16'h322A
`define CUBE_LUT_323F 16'h322B
`define CUBE_LUT_3240 16'h322C
`define CUBE_LUT_3241 16'h322D
`define CUBE_LUT_3242 16'h322E
`define CUBE_LUT_3243 16'h322F
`define CUBE_LUT_3244 16'h3230
`define CUBE_LUT_3245 16'h3231
`define CUBE_LUT_3246 16'h3232
`define CUBE_LUT_3247 16'h3233
`define CUBE_LUT_3248 16'h3234
`define CUBE_LUT_3249 16'h3235
`define CUBE_LUT_324A 16'h3236
`define CUBE_LUT_324B 16'h3237
`define CUBE_LUT_324C 16'h3238
`define CUBE_LUT_324D 16'h3238
`define CUBE_LUT_324E 16'h3239
`define CUBE_LUT_324F 16'h323A
`define CUBE_LUT_3250 16'h323B
`define CUBE_LUT_3251 16'h323C
`define CUBE_LUT_3252 16'h323D
`define CUBE_LUT_3253 16'h323E
`define CUBE_LUT_3254 16'h323F
`define CUBE_LUT_3255 16'h3240
`define CUBE_LUT_3256 16'h3241
`define CUBE_LUT_3257 16'h3242
`define CUBE_LUT_3258 16'h3243
`define CUBE_LUT_3259 16'h3244
`define CUBE_LUT_325A 16'h3245
`define CUBE_LUT_325B 16'h3246
`define CUBE_LUT_325C 16'h3247
`define CUBE_LUT_325D 16'h3248
`define CUBE_LUT_325E 16'h3249
`define CUBE_LUT_325F 16'h324A
`define CUBE_LUT_3260 16'h324B
`define CUBE_LUT_3261 16'h324C
`define CUBE_LUT_3262 16'h324D
`define CUBE_LUT_3263 16'h324E
`define CUBE_LUT_3264 16'h324F
`define CUBE_LUT_3265 16'h3250
`define CUBE_LUT_3266 16'h3251
`define CUBE_LUT_3267 16'h3251
`define CUBE_LUT_3268 16'h3252
`define CUBE_LUT_3269 16'h3253
`define CUBE_LUT_326A 16'h3254
`define CUBE_LUT_326B 16'h3255
`define CUBE_LUT_326C 16'h3256
`define CUBE_LUT_326D 16'h3257
`define CUBE_LUT_326E 16'h3258
`define CUBE_LUT_326F 16'h3259
`define CUBE_LUT_3270 16'h325A
`define CUBE_LUT_3271 16'h325B
`define CUBE_LUT_3272 16'h325C
`define CUBE_LUT_3273 16'h325D
`define CUBE_LUT_3274 16'h325E
`define CUBE_LUT_3275 16'h325F
`define CUBE_LUT_3276 16'h3260
`define CUBE_LUT_3277 16'h3261
`define CUBE_LUT_3278 16'h3262
`define CUBE_LUT_3279 16'h3263
`define CUBE_LUT_327A 16'h3264
`define CUBE_LUT_327B 16'h3265
`define CUBE_LUT_327C 16'h3266
`define CUBE_LUT_327D 16'h3267
`define CUBE_LUT_327E 16'h3268
`define CUBE_LUT_327F 16'h3269
`define CUBE_LUT_3280 16'h3269
`define CUBE_LUT_3281 16'h326A
`define CUBE_LUT_3282 16'h326B
`define CUBE_LUT_3283 16'h326C
`define CUBE_LUT_3284 16'h326D
`define CUBE_LUT_3285 16'h326E
`define CUBE_LUT_3286 16'h326F
`define CUBE_LUT_3287 16'h3270
`define CUBE_LUT_3288 16'h3271
`define CUBE_LUT_3289 16'h3272
`define CUBE_LUT_328A 16'h3273
`define CUBE_LUT_328B 16'h3274
`define CUBE_LUT_328C 16'h3275
`define CUBE_LUT_328D 16'h3276
`define CUBE_LUT_328E 16'h3277
`define CUBE_LUT_328F 16'h3278
`define CUBE_LUT_3290 16'h3279
`define CUBE_LUT_3291 16'h327A
`define CUBE_LUT_3292 16'h327B
`define CUBE_LUT_3293 16'h327C
`define CUBE_LUT_3294 16'h327D
`define CUBE_LUT_3295 16'h327E
`define CUBE_LUT_3296 16'h327F
`define CUBE_LUT_3297 16'h3280
`define CUBE_LUT_3298 16'h3281
`define CUBE_LUT_3299 16'h3281
`define CUBE_LUT_329A 16'h3282
`define CUBE_LUT_329B 16'h3283
`define CUBE_LUT_329C 16'h3284
`define CUBE_LUT_329D 16'h3285
`define CUBE_LUT_329E 16'h3286
`define CUBE_LUT_329F 16'h3287
`define CUBE_LUT_32A0 16'h3288
`define CUBE_LUT_32A1 16'h3289
`define CUBE_LUT_32A2 16'h328A
`define CUBE_LUT_32A3 16'h328B
`define CUBE_LUT_32A4 16'h328C
`define CUBE_LUT_32A5 16'h328D
`define CUBE_LUT_32A6 16'h328E
`define CUBE_LUT_32A7 16'h328F
`define CUBE_LUT_32A8 16'h3290
`define CUBE_LUT_32A9 16'h3291
`define CUBE_LUT_32AA 16'h3292
`define CUBE_LUT_32AB 16'h3293
`define CUBE_LUT_32AC 16'h3294
`define CUBE_LUT_32AD 16'h3295
`define CUBE_LUT_32AE 16'h3296
`define CUBE_LUT_32AF 16'h3297
`define CUBE_LUT_32B0 16'h3298
`define CUBE_LUT_32B1 16'h3298
`define CUBE_LUT_32B2 16'h3299
`define CUBE_LUT_32B3 16'h329A
`define CUBE_LUT_32B4 16'h329B
`define CUBE_LUT_32B5 16'h329C
`define CUBE_LUT_32B6 16'h329D
`define CUBE_LUT_32B7 16'h329E
`define CUBE_LUT_32B8 16'h329F
`define CUBE_LUT_32B9 16'h32A0
`define CUBE_LUT_32BA 16'h32A1
`define CUBE_LUT_32BB 16'h32A2
`define CUBE_LUT_32BC 16'h32A3
`define CUBE_LUT_32BD 16'h32A4
`define CUBE_LUT_32BE 16'h32A5
`define CUBE_LUT_32BF 16'h32A6
`define CUBE_LUT_32C0 16'h32A7
`define CUBE_LUT_32C1 16'h32A8
`define CUBE_LUT_32C2 16'h32A9
`define CUBE_LUT_32C3 16'h32AA
`define CUBE_LUT_32C4 16'h32AB
`define CUBE_LUT_32C5 16'h32AC
`define CUBE_LUT_32C6 16'h32AD
`define CUBE_LUT_32C7 16'h32AE
`define CUBE_LUT_32C8 16'h32AE
`define CUBE_LUT_32C9 16'h32AF
`define CUBE_LUT_32CA 16'h32B0
`define CUBE_LUT_32CB 16'h32B1
`define CUBE_LUT_32CC 16'h32B2
`define CUBE_LUT_32CD 16'h32B3
`define CUBE_LUT_32CE 16'h32B4
`define CUBE_LUT_32CF 16'h32B5
`define CUBE_LUT_32D0 16'h32B6
`define CUBE_LUT_32D1 16'h32B7
`define CUBE_LUT_32D2 16'h32B8
`define CUBE_LUT_32D3 16'h32B9
`define CUBE_LUT_32D4 16'h32BA
`define CUBE_LUT_32D5 16'h32BB
`define CUBE_LUT_32D6 16'h32BC
`define CUBE_LUT_32D7 16'h32BD
`define CUBE_LUT_32D8 16'h32BE
`define CUBE_LUT_32D9 16'h32BF
`define CUBE_LUT_32DA 16'h32C0
`define CUBE_LUT_32DB 16'h32C1
`define CUBE_LUT_32DC 16'h32C2
`define CUBE_LUT_32DD 16'h32C3
`define CUBE_LUT_32DE 16'h32C4
`define CUBE_LUT_32DF 16'h32C4
`define CUBE_LUT_32E0 16'h32C5
`define CUBE_LUT_32E1 16'h32C6
`define CUBE_LUT_32E2 16'h32C7
`define CUBE_LUT_32E3 16'h32C8
`define CUBE_LUT_32E4 16'h32C9
`define CUBE_LUT_32E5 16'h32CA
`define CUBE_LUT_32E6 16'h32CB
`define CUBE_LUT_32E7 16'h32CC
`define CUBE_LUT_32E8 16'h32CD
`define CUBE_LUT_32E9 16'h32CE
`define CUBE_LUT_32EA 16'h32CF
`define CUBE_LUT_32EB 16'h32D0
`define CUBE_LUT_32EC 16'h32D1
`define CUBE_LUT_32ED 16'h32D2
`define CUBE_LUT_32EE 16'h32D3
`define CUBE_LUT_32EF 16'h32D4
`define CUBE_LUT_32F0 16'h32D5
`define CUBE_LUT_32F1 16'h32D6
`define CUBE_LUT_32F2 16'h32D7
`define CUBE_LUT_32F3 16'h32D8
`define CUBE_LUT_32F4 16'h32D9
`define CUBE_LUT_32F5 16'h32D9
`define CUBE_LUT_32F6 16'h32DA
`define CUBE_LUT_32F7 16'h32DB
`define CUBE_LUT_32F8 16'h32DC
`define CUBE_LUT_32F9 16'h32DD
`define CUBE_LUT_32FA 16'h32DE
`define CUBE_LUT_32FB 16'h32DF
`define CUBE_LUT_32FC 16'h32E0
`define CUBE_LUT_32FD 16'h32E1
`define CUBE_LUT_32FE 16'h32E2
`define CUBE_LUT_32FF 16'h32E3
`define CUBE_LUT_3300 16'h32E4
`define CUBE_LUT_3301 16'h32E5
`define CUBE_LUT_3302 16'h32E6
`define CUBE_LUT_3303 16'h32E7
`define CUBE_LUT_3304 16'h32E8
`define CUBE_LUT_3305 16'h32E9
`define CUBE_LUT_3306 16'h32EA
`define CUBE_LUT_3307 16'h32EB
`define CUBE_LUT_3308 16'h32EC
`define CUBE_LUT_3309 16'h32ED
`define CUBE_LUT_330A 16'h32ED
`define CUBE_LUT_330B 16'h32EE
`define CUBE_LUT_330C 16'h32EF
`define CUBE_LUT_330D 16'h32F0
`define CUBE_LUT_330E 16'h32F1
`define CUBE_LUT_330F 16'h32F2
`define CUBE_LUT_3310 16'h32F3
`define CUBE_LUT_3311 16'h32F4
`define CUBE_LUT_3312 16'h32F5
`define CUBE_LUT_3313 16'h32F6
`define CUBE_LUT_3314 16'h32F7
`define CUBE_LUT_3315 16'h32F8
`define CUBE_LUT_3316 16'h32F9
`define CUBE_LUT_3317 16'h32FA
`define CUBE_LUT_3318 16'h32FB
`define CUBE_LUT_3319 16'h32FC
`define CUBE_LUT_331A 16'h32FD
`define CUBE_LUT_331B 16'h32FE
`define CUBE_LUT_331C 16'h32FF
`define CUBE_LUT_331D 16'h3300
`define CUBE_LUT_331E 16'h3301
`define CUBE_LUT_331F 16'h3301
`define CUBE_LUT_3320 16'h3302
`define CUBE_LUT_3321 16'h3303
`define CUBE_LUT_3322 16'h3304
`define CUBE_LUT_3323 16'h3305
`define CUBE_LUT_3324 16'h3306
`define CUBE_LUT_3325 16'h3307
`define CUBE_LUT_3326 16'h3308
`define CUBE_LUT_3327 16'h3309
`define CUBE_LUT_3328 16'h330A
`define CUBE_LUT_3329 16'h330B
`define CUBE_LUT_332A 16'h330C
`define CUBE_LUT_332B 16'h330D
`define CUBE_LUT_332C 16'h330E
`define CUBE_LUT_332D 16'h330F
`define CUBE_LUT_332E 16'h3310
`define CUBE_LUT_332F 16'h3311
`define CUBE_LUT_3330 16'h3312
`define CUBE_LUT_3331 16'h3313
`define CUBE_LUT_3332 16'h3314
`define CUBE_LUT_3333 16'h3315
`define CUBE_LUT_3334 16'h3315
`define CUBE_LUT_3335 16'h3316
`define CUBE_LUT_3336 16'h3317
`define CUBE_LUT_3337 16'h3318
`define CUBE_LUT_3338 16'h3319
`define CUBE_LUT_3339 16'h331A
`define CUBE_LUT_333A 16'h331B
`define CUBE_LUT_333B 16'h331C
`define CUBE_LUT_333C 16'h331D
`define CUBE_LUT_333D 16'h331E
`define CUBE_LUT_333E 16'h331F
`define CUBE_LUT_333F 16'h3320
`define CUBE_LUT_3340 16'h3321
`define CUBE_LUT_3341 16'h3322
`define CUBE_LUT_3342 16'h3323
`define CUBE_LUT_3343 16'h3324
`define CUBE_LUT_3344 16'h3325
`define CUBE_LUT_3345 16'h3326
`define CUBE_LUT_3346 16'h3327
`define CUBE_LUT_3347 16'h3328
`define CUBE_LUT_3348 16'h3328
`define CUBE_LUT_3349 16'h3329
`define CUBE_LUT_334A 16'h332A
`define CUBE_LUT_334B 16'h332B
`define CUBE_LUT_334C 16'h332C
`define CUBE_LUT_334D 16'h332D
`define CUBE_LUT_334E 16'h332E
`define CUBE_LUT_334F 16'h332F
`define CUBE_LUT_3350 16'h3330
`define CUBE_LUT_3351 16'h3331
`define CUBE_LUT_3352 16'h3332
`define CUBE_LUT_3353 16'h3333
`define CUBE_LUT_3354 16'h3334
`define CUBE_LUT_3355 16'h3335
`define CUBE_LUT_3356 16'h3336
`define CUBE_LUT_3357 16'h3337
`define CUBE_LUT_3358 16'h3338
`define CUBE_LUT_3359 16'h3339
`define CUBE_LUT_335A 16'h333A
`define CUBE_LUT_335B 16'h333B
`define CUBE_LUT_335C 16'h333B
`define CUBE_LUT_335D 16'h333C
`define CUBE_LUT_335E 16'h333D
`define CUBE_LUT_335F 16'h333E
`define CUBE_LUT_3360 16'h333F
`define CUBE_LUT_3361 16'h3340
`define CUBE_LUT_3362 16'h3341
`define CUBE_LUT_3363 16'h3342
`define CUBE_LUT_3364 16'h3343
`define CUBE_LUT_3365 16'h3344
`define CUBE_LUT_3366 16'h3345
`define CUBE_LUT_3367 16'h3346
`define CUBE_LUT_3368 16'h3347
`define CUBE_LUT_3369 16'h3348
`define CUBE_LUT_336A 16'h3349
`define CUBE_LUT_336B 16'h334A
`define CUBE_LUT_336C 16'h334B
`define CUBE_LUT_336D 16'h334C
`define CUBE_LUT_336E 16'h334D
`define CUBE_LUT_336F 16'h334D
`define CUBE_LUT_3370 16'h334E
`define CUBE_LUT_3371 16'h334F
`define CUBE_LUT_3372 16'h3350
`define CUBE_LUT_3373 16'h3351
`define CUBE_LUT_3374 16'h3352
`define CUBE_LUT_3375 16'h3353
`define CUBE_LUT_3376 16'h3354
`define CUBE_LUT_3377 16'h3355
`define CUBE_LUT_3378 16'h3356
`define CUBE_LUT_3379 16'h3357
`define CUBE_LUT_337A 16'h3358
`define CUBE_LUT_337B 16'h3359
`define CUBE_LUT_337C 16'h335A
`define CUBE_LUT_337D 16'h335B
`define CUBE_LUT_337E 16'h335C
`define CUBE_LUT_337F 16'h335D
`define CUBE_LUT_3380 16'h335E
`define CUBE_LUT_3381 16'h335F
`define CUBE_LUT_3382 16'h335F
`define CUBE_LUT_3383 16'h3360
`define CUBE_LUT_3384 16'h3361
`define CUBE_LUT_3385 16'h3362
`define CUBE_LUT_3386 16'h3363
`define CUBE_LUT_3387 16'h3364
`define CUBE_LUT_3388 16'h3365
`define CUBE_LUT_3389 16'h3366
`define CUBE_LUT_338A 16'h3367
`define CUBE_LUT_338B 16'h3368
`define CUBE_LUT_338C 16'h3369
`define CUBE_LUT_338D 16'h336A
`define CUBE_LUT_338E 16'h336B
`define CUBE_LUT_338F 16'h336C
`define CUBE_LUT_3390 16'h336D
`define CUBE_LUT_3391 16'h336E
`define CUBE_LUT_3392 16'h336F
`define CUBE_LUT_3393 16'h3370
`define CUBE_LUT_3394 16'h3371
`define CUBE_LUT_3395 16'h3371
`define CUBE_LUT_3396 16'h3372
`define CUBE_LUT_3397 16'h3373
`define CUBE_LUT_3398 16'h3374
`define CUBE_LUT_3399 16'h3375
`define CUBE_LUT_339A 16'h3376
`define CUBE_LUT_339B 16'h3377
`define CUBE_LUT_339C 16'h3378
`define CUBE_LUT_339D 16'h3379
`define CUBE_LUT_339E 16'h337A
`define CUBE_LUT_339F 16'h337B
`define CUBE_LUT_33A0 16'h337C
`define CUBE_LUT_33A1 16'h337D
`define CUBE_LUT_33A2 16'h337E
`define CUBE_LUT_33A3 16'h337F
`define CUBE_LUT_33A4 16'h3380
`define CUBE_LUT_33A5 16'h3381
`define CUBE_LUT_33A6 16'h3382
`define CUBE_LUT_33A7 16'h3382
`define CUBE_LUT_33A8 16'h3383
`define CUBE_LUT_33A9 16'h3384
`define CUBE_LUT_33AA 16'h3385
`define CUBE_LUT_33AB 16'h3386
`define CUBE_LUT_33AC 16'h3387
`define CUBE_LUT_33AD 16'h3388
`define CUBE_LUT_33AE 16'h3389
`define CUBE_LUT_33AF 16'h338A
`define CUBE_LUT_33B0 16'h338B
`define CUBE_LUT_33B1 16'h338C
`define CUBE_LUT_33B2 16'h338D
`define CUBE_LUT_33B3 16'h338E
`define CUBE_LUT_33B4 16'h338F
`define CUBE_LUT_33B5 16'h3390
`define CUBE_LUT_33B6 16'h3391
`define CUBE_LUT_33B7 16'h3392
`define CUBE_LUT_33B8 16'h3393
`define CUBE_LUT_33B9 16'h3393
`define CUBE_LUT_33BA 16'h3394
`define CUBE_LUT_33BB 16'h3395
`define CUBE_LUT_33BC 16'h3396
`define CUBE_LUT_33BD 16'h3397
`define CUBE_LUT_33BE 16'h3398
`define CUBE_LUT_33BF 16'h3399
`define CUBE_LUT_33C0 16'h339A
`define CUBE_LUT_33C1 16'h339B
`define CUBE_LUT_33C2 16'h339C
`define CUBE_LUT_33C3 16'h339D
`define CUBE_LUT_33C4 16'h339E
`define CUBE_LUT_33C5 16'h339F
`define CUBE_LUT_33C6 16'h33A0
`define CUBE_LUT_33C7 16'h33A1
`define CUBE_LUT_33C8 16'h33A2
`define CUBE_LUT_33C9 16'h33A3
`define CUBE_LUT_33CA 16'h33A4
`define CUBE_LUT_33CB 16'h33A4
`define CUBE_LUT_33CC 16'h33A5
`define CUBE_LUT_33CD 16'h33A6
`define CUBE_LUT_33CE 16'h33A7
`define CUBE_LUT_33CF 16'h33A8
`define CUBE_LUT_33D0 16'h33A9
`define CUBE_LUT_33D1 16'h33AA
`define CUBE_LUT_33D2 16'h33AB
`define CUBE_LUT_33D3 16'h33AC
`define CUBE_LUT_33D4 16'h33AD
`define CUBE_LUT_33D5 16'h33AE
`define CUBE_LUT_33D6 16'h33AF
`define CUBE_LUT_33D7 16'h33B0
`define CUBE_LUT_33D8 16'h33B1
`define CUBE_LUT_33D9 16'h33B2
`define CUBE_LUT_33DA 16'h33B3
`define CUBE_LUT_33DB 16'h33B4
`define CUBE_LUT_33DC 16'h33B4
`define CUBE_LUT_33DD 16'h33B5
`define CUBE_LUT_33DE 16'h33B6
`define CUBE_LUT_33DF 16'h33B7
`define CUBE_LUT_33E0 16'h33B8
`define CUBE_LUT_33E1 16'h33B9
`define CUBE_LUT_33E2 16'h33BA
`define CUBE_LUT_33E3 16'h33BB
`define CUBE_LUT_33E4 16'h33BC
`define CUBE_LUT_33E5 16'h33BD
`define CUBE_LUT_33E6 16'h33BE
`define CUBE_LUT_33E7 16'h33BF
`define CUBE_LUT_33E8 16'h33C0
`define CUBE_LUT_33E9 16'h33C1
`define CUBE_LUT_33EA 16'h33C2
`define CUBE_LUT_33EB 16'h33C3
`define CUBE_LUT_33EC 16'h33C4
`define CUBE_LUT_33ED 16'h33C5
`define CUBE_LUT_33EE 16'h33C5
`define CUBE_LUT_33EF 16'h33C6
`define CUBE_LUT_33F0 16'h33C7
`define CUBE_LUT_33F1 16'h33C8
`define CUBE_LUT_33F2 16'h33C9
`define CUBE_LUT_33F3 16'h33CA
`define CUBE_LUT_33F4 16'h33CB
`define CUBE_LUT_33F5 16'h33CC
`define CUBE_LUT_33F6 16'h33CD
`define CUBE_LUT_33F7 16'h33CE
`define CUBE_LUT_33F8 16'h33CF
`define CUBE_LUT_33F9 16'h33D0
`define CUBE_LUT_33FA 16'h33D1
`define CUBE_LUT_33FB 16'h33D2
`define CUBE_LUT_33FC 16'h33D3
`define CUBE_LUT_33FD 16'h33D4
`define CUBE_LUT_33FE 16'h33D4
`define CUBE_LUT_33FF 16'h33D5
`define CUBE_LUT_3400 16'h33D6
`define CUBE_LUT_3401 16'h33D8
`define CUBE_LUT_3402 16'h33DA
`define CUBE_LUT_3403 16'h33DC
`define CUBE_LUT_3404 16'h33DE
`define CUBE_LUT_3405 16'h33E0
`define CUBE_LUT_3406 16'h33E2
`define CUBE_LUT_3407 16'h33E4
`define CUBE_LUT_3408 16'h33E5
`define CUBE_LUT_3409 16'h33E7
`define CUBE_LUT_340A 16'h33E9
`define CUBE_LUT_340B 16'h33EB
`define CUBE_LUT_340C 16'h33ED
`define CUBE_LUT_340D 16'h33EF
`define CUBE_LUT_340E 16'h33F1
`define CUBE_LUT_340F 16'h33F3
`define CUBE_LUT_3410 16'h33F4
`define CUBE_LUT_3411 16'h33F6
`define CUBE_LUT_3412 16'h33F8
`define CUBE_LUT_3413 16'h33FA
`define CUBE_LUT_3414 16'h33FC
`define CUBE_LUT_3415 16'h33FE
`define CUBE_LUT_3416 16'h3400
`define CUBE_LUT_3417 16'h3401
`define CUBE_LUT_3418 16'h3402
`define CUBE_LUT_3419 16'h3403
`define CUBE_LUT_341A 16'h3404
`define CUBE_LUT_341B 16'h3405
`define CUBE_LUT_341C 16'h3405
`define CUBE_LUT_341D 16'h3406
`define CUBE_LUT_341E 16'h3407
`define CUBE_LUT_341F 16'h3408
`define CUBE_LUT_3420 16'h3409
`define CUBE_LUT_3421 16'h340A
`define CUBE_LUT_3422 16'h340B
`define CUBE_LUT_3423 16'h340C
`define CUBE_LUT_3424 16'h340D
`define CUBE_LUT_3425 16'h340E
`define CUBE_LUT_3426 16'h340F
`define CUBE_LUT_3427 16'h3410
`define CUBE_LUT_3428 16'h3411
`define CUBE_LUT_3429 16'h3412
`define CUBE_LUT_342A 16'h3413
`define CUBE_LUT_342B 16'h3414
`define CUBE_LUT_342C 16'h3414
`define CUBE_LUT_342D 16'h3415
`define CUBE_LUT_342E 16'h3416
`define CUBE_LUT_342F 16'h3417
`define CUBE_LUT_3430 16'h3418
`define CUBE_LUT_3431 16'h3419
`define CUBE_LUT_3432 16'h341A
`define CUBE_LUT_3433 16'h341B
`define CUBE_LUT_3434 16'h341C
`define CUBE_LUT_3435 16'h341D
`define CUBE_LUT_3436 16'h341E
`define CUBE_LUT_3437 16'h341F
`define CUBE_LUT_3438 16'h3420
`define CUBE_LUT_3439 16'h3421
`define CUBE_LUT_343A 16'h3422
`define CUBE_LUT_343B 16'h3422
`define CUBE_LUT_343C 16'h3423
`define CUBE_LUT_343D 16'h3424
`define CUBE_LUT_343E 16'h3425
`define CUBE_LUT_343F 16'h3426
`define CUBE_LUT_3440 16'h3427
`define CUBE_LUT_3441 16'h3428
`define CUBE_LUT_3442 16'h3429
`define CUBE_LUT_3443 16'h342A
`define CUBE_LUT_3444 16'h342B
`define CUBE_LUT_3445 16'h342C
`define CUBE_LUT_3446 16'h342D
`define CUBE_LUT_3447 16'h342E
`define CUBE_LUT_3448 16'h342F
`define CUBE_LUT_3449 16'h3430
`define CUBE_LUT_344A 16'h3430
`define CUBE_LUT_344B 16'h3431
`define CUBE_LUT_344C 16'h3432
`define CUBE_LUT_344D 16'h3433
`define CUBE_LUT_344E 16'h3434
`define CUBE_LUT_344F 16'h3435
`define CUBE_LUT_3450 16'h3436
`define CUBE_LUT_3451 16'h3437
`define CUBE_LUT_3452 16'h3438
`define CUBE_LUT_3453 16'h3439
`define CUBE_LUT_3454 16'h343A
`define CUBE_LUT_3455 16'h343B
`define CUBE_LUT_3456 16'h343C
`define CUBE_LUT_3457 16'h343D
`define CUBE_LUT_3458 16'h343D
`define CUBE_LUT_3459 16'h343E
`define CUBE_LUT_345A 16'h343F
`define CUBE_LUT_345B 16'h3440
`define CUBE_LUT_345C 16'h3441
`define CUBE_LUT_345D 16'h3442
`define CUBE_LUT_345E 16'h3443
`define CUBE_LUT_345F 16'h3444
`define CUBE_LUT_3460 16'h3445
`define CUBE_LUT_3461 16'h3446
`define CUBE_LUT_3462 16'h3447
`define CUBE_LUT_3463 16'h3448
`define CUBE_LUT_3464 16'h3449
`define CUBE_LUT_3465 16'h344A
`define CUBE_LUT_3466 16'h344A
`define CUBE_LUT_3467 16'h344B
`define CUBE_LUT_3468 16'h344C
`define CUBE_LUT_3469 16'h344D
`define CUBE_LUT_346A 16'h344E
`define CUBE_LUT_346B 16'h344F
`define CUBE_LUT_346C 16'h3450
`define CUBE_LUT_346D 16'h3451
`define CUBE_LUT_346E 16'h3452
`define CUBE_LUT_346F 16'h3453
`define CUBE_LUT_3470 16'h3454
`define CUBE_LUT_3471 16'h3455
`define CUBE_LUT_3472 16'h3456
`define CUBE_LUT_3473 16'h3457
`define CUBE_LUT_3474 16'h3457
`define CUBE_LUT_3475 16'h3458
`define CUBE_LUT_3476 16'h3459
`define CUBE_LUT_3477 16'h345A
`define CUBE_LUT_3478 16'h345B
`define CUBE_LUT_3479 16'h345C
`define CUBE_LUT_347A 16'h345D
`define CUBE_LUT_347B 16'h345E
`define CUBE_LUT_347C 16'h345F
`define CUBE_LUT_347D 16'h3460
`define CUBE_LUT_347E 16'h3461
`define CUBE_LUT_347F 16'h3462
`define CUBE_LUT_3480 16'h3463
`define CUBE_LUT_3481 16'h3463
`define CUBE_LUT_3482 16'h3464
`define CUBE_LUT_3483 16'h3465
`define CUBE_LUT_3484 16'h3466
`define CUBE_LUT_3485 16'h3467
`define CUBE_LUT_3486 16'h3468
`define CUBE_LUT_3487 16'h3469
`define CUBE_LUT_3488 16'h346A
`define CUBE_LUT_3489 16'h346B
`define CUBE_LUT_348A 16'h346C
`define CUBE_LUT_348B 16'h346D
`define CUBE_LUT_348C 16'h346E
`define CUBE_LUT_348D 16'h346F
`define CUBE_LUT_348E 16'h346F
`define CUBE_LUT_348F 16'h3470
`define CUBE_LUT_3490 16'h3471
`define CUBE_LUT_3491 16'h3472
`define CUBE_LUT_3492 16'h3473
`define CUBE_LUT_3493 16'h3474
`define CUBE_LUT_3494 16'h3475
`define CUBE_LUT_3495 16'h3476
`define CUBE_LUT_3496 16'h3477
`define CUBE_LUT_3497 16'h3478
`define CUBE_LUT_3498 16'h3479
`define CUBE_LUT_3499 16'h347A
`define CUBE_LUT_349A 16'h347B
`define CUBE_LUT_349B 16'h347B
`define CUBE_LUT_349C 16'h347C
`define CUBE_LUT_349D 16'h347D
`define CUBE_LUT_349E 16'h347E
`define CUBE_LUT_349F 16'h347F
`define CUBE_LUT_34A0 16'h3480
`define CUBE_LUT_34A1 16'h3481
`define CUBE_LUT_34A2 16'h3482
`define CUBE_LUT_34A3 16'h3483
`define CUBE_LUT_34A4 16'h3484
`define CUBE_LUT_34A5 16'h3485
`define CUBE_LUT_34A6 16'h3486
`define CUBE_LUT_34A7 16'h3487
`define CUBE_LUT_34A8 16'h3487
`define CUBE_LUT_34A9 16'h3488
`define CUBE_LUT_34AA 16'h3489
`define CUBE_LUT_34AB 16'h348A
`define CUBE_LUT_34AC 16'h348B
`define CUBE_LUT_34AD 16'h348C
`define CUBE_LUT_34AE 16'h348D
`define CUBE_LUT_34AF 16'h348E
`define CUBE_LUT_34B0 16'h348F
`define CUBE_LUT_34B1 16'h3490
`define CUBE_LUT_34B2 16'h3491
`define CUBE_LUT_34B3 16'h3492
`define CUBE_LUT_34B4 16'h3492
`define CUBE_LUT_34B5 16'h3493
`define CUBE_LUT_34B6 16'h3494
`define CUBE_LUT_34B7 16'h3495
`define CUBE_LUT_34B8 16'h3496
`define CUBE_LUT_34B9 16'h3497
`define CUBE_LUT_34BA 16'h3498
`define CUBE_LUT_34BB 16'h3499
`define CUBE_LUT_34BC 16'h349A
`define CUBE_LUT_34BD 16'h349B
`define CUBE_LUT_34BE 16'h349C
`define CUBE_LUT_34BF 16'h349D
`define CUBE_LUT_34C0 16'h349D
`define CUBE_LUT_34C1 16'h349E
`define CUBE_LUT_34C2 16'h349F
`define CUBE_LUT_34C3 16'h34A0
`define CUBE_LUT_34C4 16'h34A1
`define CUBE_LUT_34C5 16'h34A2
`define CUBE_LUT_34C6 16'h34A3
`define CUBE_LUT_34C7 16'h34A4
`define CUBE_LUT_34C8 16'h34A5
`define CUBE_LUT_34C9 16'h34A6
`define CUBE_LUT_34CA 16'h34A7
`define CUBE_LUT_34CB 16'h34A8
`define CUBE_LUT_34CC 16'h34A8
`define CUBE_LUT_34CD 16'h34A9
`define CUBE_LUT_34CE 16'h34AA
`define CUBE_LUT_34CF 16'h34AB
`define CUBE_LUT_34D0 16'h34AC
`define CUBE_LUT_34D1 16'h34AD
`define CUBE_LUT_34D2 16'h34AE
`define CUBE_LUT_34D3 16'h34AF
`define CUBE_LUT_34D4 16'h34B0
`define CUBE_LUT_34D5 16'h34B1
`define CUBE_LUT_34D6 16'h34B2
`define CUBE_LUT_34D7 16'h34B3
`define CUBE_LUT_34D8 16'h34B3
`define CUBE_LUT_34D9 16'h34B4
`define CUBE_LUT_34DA 16'h34B5
`define CUBE_LUT_34DB 16'h34B6
`define CUBE_LUT_34DC 16'h34B7
`define CUBE_LUT_34DD 16'h34B8
`define CUBE_LUT_34DE 16'h34B9
`define CUBE_LUT_34DF 16'h34BA
`define CUBE_LUT_34E0 16'h34BB
`define CUBE_LUT_34E1 16'h34BC
`define CUBE_LUT_34E2 16'h34BD
`define CUBE_LUT_34E3 16'h34BE
`define CUBE_LUT_34E4 16'h34BE
`define CUBE_LUT_34E5 16'h34BF
`define CUBE_LUT_34E6 16'h34C0
`define CUBE_LUT_34E7 16'h34C1
`define CUBE_LUT_34E8 16'h34C2
`define CUBE_LUT_34E9 16'h34C3
`define CUBE_LUT_34EA 16'h34C4
`define CUBE_LUT_34EB 16'h34C5
`define CUBE_LUT_34EC 16'h34C6
`define CUBE_LUT_34ED 16'h34C7
`define CUBE_LUT_34EE 16'h34C8
`define CUBE_LUT_34EF 16'h34C8
`define CUBE_LUT_34F0 16'h34C9
`define CUBE_LUT_34F1 16'h34CA
`define CUBE_LUT_34F2 16'h34CB
`define CUBE_LUT_34F3 16'h34CC
`define CUBE_LUT_34F4 16'h34CD
`define CUBE_LUT_34F5 16'h34CE
`define CUBE_LUT_34F6 16'h34CF
`define CUBE_LUT_34F7 16'h34D0
`define CUBE_LUT_34F8 16'h34D1
`define CUBE_LUT_34F9 16'h34D2
`define CUBE_LUT_34FA 16'h34D2
`define CUBE_LUT_34FB 16'h34D3
`define CUBE_LUT_34FC 16'h34D4
`define CUBE_LUT_34FD 16'h34D5
`define CUBE_LUT_34FE 16'h34D6
`define CUBE_LUT_34FF 16'h34D7
`define CUBE_LUT_3500 16'h34D8
`define CUBE_LUT_3501 16'h34D9
`define CUBE_LUT_3502 16'h34DA
`define CUBE_LUT_3503 16'h34DB
`define CUBE_LUT_3504 16'h34DC
`define CUBE_LUT_3505 16'h34DC
`define CUBE_LUT_3506 16'h34DD
`define CUBE_LUT_3507 16'h34DE
`define CUBE_LUT_3508 16'h34DF
`define CUBE_LUT_3509 16'h34E0
`define CUBE_LUT_350A 16'h34E1
`define CUBE_LUT_350B 16'h34E2
`define CUBE_LUT_350C 16'h34E3
`define CUBE_LUT_350D 16'h34E4
`define CUBE_LUT_350E 16'h34E5
`define CUBE_LUT_350F 16'h34E6
`define CUBE_LUT_3510 16'h34E6
`define CUBE_LUT_3511 16'h34E7
`define CUBE_LUT_3512 16'h34E8
`define CUBE_LUT_3513 16'h34E9
`define CUBE_LUT_3514 16'h34EA
`define CUBE_LUT_3515 16'h34EB
`define CUBE_LUT_3516 16'h34EC
`define CUBE_LUT_3517 16'h34ED
`define CUBE_LUT_3518 16'h34EE
`define CUBE_LUT_3519 16'h34EF
`define CUBE_LUT_351A 16'h34EF
`define CUBE_LUT_351B 16'h34F0
`define CUBE_LUT_351C 16'h34F1
`define CUBE_LUT_351D 16'h34F2
`define CUBE_LUT_351E 16'h34F3
`define CUBE_LUT_351F 16'h34F4
`define CUBE_LUT_3520 16'h34F5
`define CUBE_LUT_3521 16'h34F6
`define CUBE_LUT_3522 16'h34F7
`define CUBE_LUT_3523 16'h34F8
`define CUBE_LUT_3524 16'h34F9
`define CUBE_LUT_3525 16'h34F9
`define CUBE_LUT_3526 16'h34FA
`define CUBE_LUT_3527 16'h34FB
`define CUBE_LUT_3528 16'h34FC
`define CUBE_LUT_3529 16'h34FD
`define CUBE_LUT_352A 16'h34FE
`define CUBE_LUT_352B 16'h34FF
`define CUBE_LUT_352C 16'h3500
`define CUBE_LUT_352D 16'h3501
`define CUBE_LUT_352E 16'h3502
`define CUBE_LUT_352F 16'h3502
`define CUBE_LUT_3530 16'h3503
`define CUBE_LUT_3531 16'h3504
`define CUBE_LUT_3532 16'h3505
`define CUBE_LUT_3533 16'h3506
`define CUBE_LUT_3534 16'h3507
`define CUBE_LUT_3535 16'h3508
`define CUBE_LUT_3536 16'h3509
`define CUBE_LUT_3537 16'h350A
`define CUBE_LUT_3538 16'h350B
`define CUBE_LUT_3539 16'h350B
`define CUBE_LUT_353A 16'h350C
`define CUBE_LUT_353B 16'h350D
`define CUBE_LUT_353C 16'h350E
`define CUBE_LUT_353D 16'h350F
`define CUBE_LUT_353E 16'h3510
`define CUBE_LUT_353F 16'h3511
`define CUBE_LUT_3540 16'h3512
`define CUBE_LUT_3541 16'h3513
`define CUBE_LUT_3542 16'h3514
`define CUBE_LUT_3543 16'h3514
`define CUBE_LUT_3544 16'h3515
`define CUBE_LUT_3545 16'h3516
`define CUBE_LUT_3546 16'h3517
`define CUBE_LUT_3547 16'h3518
`define CUBE_LUT_3548 16'h3519
`define CUBE_LUT_3549 16'h351A
`define CUBE_LUT_354A 16'h351B
`define CUBE_LUT_354B 16'h351C
`define CUBE_LUT_354C 16'h351D
`define CUBE_LUT_354D 16'h351D
`define CUBE_LUT_354E 16'h351E
`define CUBE_LUT_354F 16'h351F
`define CUBE_LUT_3550 16'h3520
`define CUBE_LUT_3551 16'h3521
`define CUBE_LUT_3552 16'h3522
`define CUBE_LUT_3553 16'h3523
`define CUBE_LUT_3554 16'h3524
`define CUBE_LUT_3555 16'h3525
`define CUBE_LUT_3556 16'h3526
`define CUBE_LUT_3557 16'h3526
`define CUBE_LUT_3558 16'h3527
`define CUBE_LUT_3559 16'h3528
`define CUBE_LUT_355A 16'h3529
`define CUBE_LUT_355B 16'h352A
`define CUBE_LUT_355C 16'h352B
`define CUBE_LUT_355D 16'h352C
`define CUBE_LUT_355E 16'h352D
`define CUBE_LUT_355F 16'h352E
`define CUBE_LUT_3560 16'h352E
`define CUBE_LUT_3561 16'h352F
`define CUBE_LUT_3562 16'h3530
`define CUBE_LUT_3563 16'h3531
`define CUBE_LUT_3564 16'h3532
`define CUBE_LUT_3565 16'h3533
`define CUBE_LUT_3566 16'h3534
`define CUBE_LUT_3567 16'h3535
`define CUBE_LUT_3568 16'h3536
`define CUBE_LUT_3569 16'h3537
`define CUBE_LUT_356A 16'h3537
`define CUBE_LUT_356B 16'h3538
`define CUBE_LUT_356C 16'h3539
`define CUBE_LUT_356D 16'h353A
`define CUBE_LUT_356E 16'h353B
`define CUBE_LUT_356F 16'h353C
`define CUBE_LUT_3570 16'h353D
`define CUBE_LUT_3571 16'h353E
`define CUBE_LUT_3572 16'h353F
`define CUBE_LUT_3573 16'h353F
`define CUBE_LUT_3574 16'h3540
`define CUBE_LUT_3575 16'h3541
`define CUBE_LUT_3576 16'h3542
`define CUBE_LUT_3577 16'h3543
`define CUBE_LUT_3578 16'h3544
`define CUBE_LUT_3579 16'h3545
`define CUBE_LUT_357A 16'h3546
`define CUBE_LUT_357B 16'h3547
`define CUBE_LUT_357C 16'h3547
`define CUBE_LUT_357D 16'h3548
`define CUBE_LUT_357E 16'h3549
`define CUBE_LUT_357F 16'h354A
`define CUBE_LUT_3580 16'h354B
`define CUBE_LUT_3581 16'h354C
`define CUBE_LUT_3582 16'h354D
`define CUBE_LUT_3583 16'h354E
`define CUBE_LUT_3584 16'h354F
`define CUBE_LUT_3585 16'h354F
`define CUBE_LUT_3586 16'h3550
`define CUBE_LUT_3587 16'h3551
`define CUBE_LUT_3588 16'h3552
`define CUBE_LUT_3589 16'h3553
`define CUBE_LUT_358A 16'h3554
`define CUBE_LUT_358B 16'h3555
`define CUBE_LUT_358C 16'h3556
`define CUBE_LUT_358D 16'h3557
`define CUBE_LUT_358E 16'h3557
`define CUBE_LUT_358F 16'h3558
`define CUBE_LUT_3590 16'h3559
`define CUBE_LUT_3591 16'h355A
`define CUBE_LUT_3592 16'h355B
`define CUBE_LUT_3593 16'h355C
`define CUBE_LUT_3594 16'h355D
`define CUBE_LUT_3595 16'h355E
`define CUBE_LUT_3596 16'h355F
`define CUBE_LUT_3597 16'h355F
`define CUBE_LUT_3598 16'h3560
`define CUBE_LUT_3599 16'h3561
`define CUBE_LUT_359A 16'h3562
`define CUBE_LUT_359B 16'h3563
`define CUBE_LUT_359C 16'h3564
`define CUBE_LUT_359D 16'h3565
`define CUBE_LUT_359E 16'h3566
`define CUBE_LUT_359F 16'h3567
`define CUBE_LUT_35A0 16'h3567
`define CUBE_LUT_35A1 16'h3568
`define CUBE_LUT_35A2 16'h3569
`define CUBE_LUT_35A3 16'h356A
`define CUBE_LUT_35A4 16'h356B
`define CUBE_LUT_35A5 16'h356C
`define CUBE_LUT_35A6 16'h356D
`define CUBE_LUT_35A7 16'h356E
`define CUBE_LUT_35A8 16'h356F
`define CUBE_LUT_35A9 16'h356F
`define CUBE_LUT_35AA 16'h3570
`define CUBE_LUT_35AB 16'h3571
`define CUBE_LUT_35AC 16'h3572
`define CUBE_LUT_35AD 16'h3573
`define CUBE_LUT_35AE 16'h3574
`define CUBE_LUT_35AF 16'h3575
`define CUBE_LUT_35B0 16'h3576
`define CUBE_LUT_35B1 16'h3577
`define CUBE_LUT_35B2 16'h3577
`define CUBE_LUT_35B3 16'h3578
`define CUBE_LUT_35B4 16'h3579
`define CUBE_LUT_35B5 16'h357A
`define CUBE_LUT_35B6 16'h357B
`define CUBE_LUT_35B7 16'h357C
`define CUBE_LUT_35B8 16'h357D
`define CUBE_LUT_35B9 16'h357E
`define CUBE_LUT_35BA 16'h357E
`define CUBE_LUT_35BB 16'h357F
`define CUBE_LUT_35BC 16'h3580
`define CUBE_LUT_35BD 16'h3581
`define CUBE_LUT_35BE 16'h3582
`define CUBE_LUT_35BF 16'h3583
`define CUBE_LUT_35C0 16'h3584
`define CUBE_LUT_35C1 16'h3585
`define CUBE_LUT_35C2 16'h3586
`define CUBE_LUT_35C3 16'h3586
`define CUBE_LUT_35C4 16'h3587
`define CUBE_LUT_35C5 16'h3588
`define CUBE_LUT_35C6 16'h3589
`define CUBE_LUT_35C7 16'h358A
`define CUBE_LUT_35C8 16'h358B
`define CUBE_LUT_35C9 16'h358C
`define CUBE_LUT_35CA 16'h358D
`define CUBE_LUT_35CB 16'h358D
`define CUBE_LUT_35CC 16'h358E
`define CUBE_LUT_35CD 16'h358F
`define CUBE_LUT_35CE 16'h3590
`define CUBE_LUT_35CF 16'h3591
`define CUBE_LUT_35D0 16'h3592
`define CUBE_LUT_35D1 16'h3593
`define CUBE_LUT_35D2 16'h3594
`define CUBE_LUT_35D3 16'h3594
`define CUBE_LUT_35D4 16'h3595
`define CUBE_LUT_35D5 16'h3596
`define CUBE_LUT_35D6 16'h3597
`define CUBE_LUT_35D7 16'h3598
`define CUBE_LUT_35D8 16'h3599
`define CUBE_LUT_35D9 16'h359A
`define CUBE_LUT_35DA 16'h359B
`define CUBE_LUT_35DB 16'h359B
`define CUBE_LUT_35DC 16'h359C
`define CUBE_LUT_35DD 16'h359D
`define CUBE_LUT_35DE 16'h359E
`define CUBE_LUT_35DF 16'h359F
`define CUBE_LUT_35E0 16'h35A0
`define CUBE_LUT_35E1 16'h35A1
`define CUBE_LUT_35E2 16'h35A2
`define CUBE_LUT_35E3 16'h35A2
`define CUBE_LUT_35E4 16'h35A3
`define CUBE_LUT_35E5 16'h35A4
`define CUBE_LUT_35E6 16'h35A5
`define CUBE_LUT_35E7 16'h35A6
`define CUBE_LUT_35E8 16'h35A7
`define CUBE_LUT_35E9 16'h35A8
`define CUBE_LUT_35EA 16'h35A9
`define CUBE_LUT_35EB 16'h35A9
`define CUBE_LUT_35EC 16'h35AA
`define CUBE_LUT_35ED 16'h35AB
`define CUBE_LUT_35EE 16'h35AC
`define CUBE_LUT_35EF 16'h35AD
`define CUBE_LUT_35F0 16'h35AE
`define CUBE_LUT_35F1 16'h35AF
`define CUBE_LUT_35F2 16'h35B0
`define CUBE_LUT_35F3 16'h35B0
`define CUBE_LUT_35F4 16'h35B1
`define CUBE_LUT_35F5 16'h35B2
`define CUBE_LUT_35F6 16'h35B3
`define CUBE_LUT_35F7 16'h35B4
`define CUBE_LUT_35F8 16'h35B5
`define CUBE_LUT_35F9 16'h35B6
`define CUBE_LUT_35FA 16'h35B7
`define CUBE_LUT_35FB 16'h35B7
`define CUBE_LUT_35FC 16'h35B8
`define CUBE_LUT_35FD 16'h35B9
`define CUBE_LUT_35FE 16'h35BA
`define CUBE_LUT_35FF 16'h35BB
`define CUBE_LUT_3600 16'h35BC
`define CUBE_LUT_3601 16'h35BD
`define CUBE_LUT_3602 16'h35BE
`define CUBE_LUT_3603 16'h35BE
`define CUBE_LUT_3604 16'h35BF
`define CUBE_LUT_3605 16'h35C0
`define CUBE_LUT_3606 16'h35C1
`define CUBE_LUT_3607 16'h35C2
`define CUBE_LUT_3608 16'h35C3
`define CUBE_LUT_3609 16'h35C4
`define CUBE_LUT_360A 16'h35C5
`define CUBE_LUT_360B 16'h35C5
`define CUBE_LUT_360C 16'h35C6
`define CUBE_LUT_360D 16'h35C7
`define CUBE_LUT_360E 16'h35C8
`define CUBE_LUT_360F 16'h35C9
`define CUBE_LUT_3610 16'h35CA
`define CUBE_LUT_3611 16'h35CB
`define CUBE_LUT_3612 16'h35CB
`define CUBE_LUT_3613 16'h35CC
`define CUBE_LUT_3614 16'h35CD
`define CUBE_LUT_3615 16'h35CE
`define CUBE_LUT_3616 16'h35CF
`define CUBE_LUT_3617 16'h35D0
`define CUBE_LUT_3618 16'h35D1
`define CUBE_LUT_3619 16'h35D2
`define CUBE_LUT_361A 16'h35D2
`define CUBE_LUT_361B 16'h35D3
`define CUBE_LUT_361C 16'h35D4
`define CUBE_LUT_361D 16'h35D5
`define CUBE_LUT_361E 16'h35D6
`define CUBE_LUT_361F 16'h35D7
`define CUBE_LUT_3620 16'h35D8
`define CUBE_LUT_3621 16'h35D9
`define CUBE_LUT_3622 16'h35D9
`define CUBE_LUT_3623 16'h35DA
`define CUBE_LUT_3624 16'h35DB
`define CUBE_LUT_3625 16'h35DC
`define CUBE_LUT_3626 16'h35DD
`define CUBE_LUT_3627 16'h35DE
`define CUBE_LUT_3628 16'h35DF
`define CUBE_LUT_3629 16'h35DF
`define CUBE_LUT_362A 16'h35E0
`define CUBE_LUT_362B 16'h35E1
`define CUBE_LUT_362C 16'h35E2
`define CUBE_LUT_362D 16'h35E3
`define CUBE_LUT_362E 16'h35E4
`define CUBE_LUT_362F 16'h35E5
`define CUBE_LUT_3630 16'h35E5
`define CUBE_LUT_3631 16'h35E6
`define CUBE_LUT_3632 16'h35E7
`define CUBE_LUT_3633 16'h35E8
`define CUBE_LUT_3634 16'h35E9
`define CUBE_LUT_3635 16'h35EA
`define CUBE_LUT_3636 16'h35EB
`define CUBE_LUT_3637 16'h35EC
`define CUBE_LUT_3638 16'h35EC
`define CUBE_LUT_3639 16'h35ED
`define CUBE_LUT_363A 16'h35EE
`define CUBE_LUT_363B 16'h35EF
`define CUBE_LUT_363C 16'h35F0
`define CUBE_LUT_363D 16'h35F1
`define CUBE_LUT_363E 16'h35F2
`define CUBE_LUT_363F 16'h35F2
`define CUBE_LUT_3640 16'h35F3
`define CUBE_LUT_3641 16'h35F4
`define CUBE_LUT_3642 16'h35F5
`define CUBE_LUT_3643 16'h35F6
`define CUBE_LUT_3644 16'h35F7
`define CUBE_LUT_3645 16'h35F8
`define CUBE_LUT_3646 16'h35F8
`define CUBE_LUT_3647 16'h35F9
`define CUBE_LUT_3648 16'h35FA
`define CUBE_LUT_3649 16'h35FB
`define CUBE_LUT_364A 16'h35FC
`define CUBE_LUT_364B 16'h35FD
`define CUBE_LUT_364C 16'h35FE
`define CUBE_LUT_364D 16'h35FE
`define CUBE_LUT_364E 16'h35FF
`define CUBE_LUT_364F 16'h3600
`define CUBE_LUT_3650 16'h3601
`define CUBE_LUT_3651 16'h3602
`define CUBE_LUT_3652 16'h3603
`define CUBE_LUT_3653 16'h3604
`define CUBE_LUT_3654 16'h3605
`define CUBE_LUT_3655 16'h3605
`define CUBE_LUT_3656 16'h3606
`define CUBE_LUT_3657 16'h3607
`define CUBE_LUT_3658 16'h3608
`define CUBE_LUT_3659 16'h3609
`define CUBE_LUT_365A 16'h360A
`define CUBE_LUT_365B 16'h360B
`define CUBE_LUT_365C 16'h360B
`define CUBE_LUT_365D 16'h360C
`define CUBE_LUT_365E 16'h360D
`define CUBE_LUT_365F 16'h360E
`define CUBE_LUT_3660 16'h360F
`define CUBE_LUT_3661 16'h3610
`define CUBE_LUT_3662 16'h3611
`define CUBE_LUT_3663 16'h3611
`define CUBE_LUT_3664 16'h3612
`define CUBE_LUT_3665 16'h3613
`define CUBE_LUT_3666 16'h3614
`define CUBE_LUT_3667 16'h3615
`define CUBE_LUT_3668 16'h3616
`define CUBE_LUT_3669 16'h3616
`define CUBE_LUT_366A 16'h3617
`define CUBE_LUT_366B 16'h3618
`define CUBE_LUT_366C 16'h3619
`define CUBE_LUT_366D 16'h361A
`define CUBE_LUT_366E 16'h361B
`define CUBE_LUT_366F 16'h361C
`define CUBE_LUT_3670 16'h361C
`define CUBE_LUT_3671 16'h361D
`define CUBE_LUT_3672 16'h361E
`define CUBE_LUT_3673 16'h361F
`define CUBE_LUT_3674 16'h3620
`define CUBE_LUT_3675 16'h3621
`define CUBE_LUT_3676 16'h3622
`define CUBE_LUT_3677 16'h3622
`define CUBE_LUT_3678 16'h3623
`define CUBE_LUT_3679 16'h3624
`define CUBE_LUT_367A 16'h3625
`define CUBE_LUT_367B 16'h3626
`define CUBE_LUT_367C 16'h3627
`define CUBE_LUT_367D 16'h3628
`define CUBE_LUT_367E 16'h3628
`define CUBE_LUT_367F 16'h3629
`define CUBE_LUT_3680 16'h362A
`define CUBE_LUT_3681 16'h362B
`define CUBE_LUT_3682 16'h362C
`define CUBE_LUT_3683 16'h362D
`define CUBE_LUT_3684 16'h362E
`define CUBE_LUT_3685 16'h362E
`define CUBE_LUT_3686 16'h362F
`define CUBE_LUT_3687 16'h3630
`define CUBE_LUT_3688 16'h3631
`define CUBE_LUT_3689 16'h3632
`define CUBE_LUT_368A 16'h3633
`define CUBE_LUT_368B 16'h3633
`define CUBE_LUT_368C 16'h3634
`define CUBE_LUT_368D 16'h3635
`define CUBE_LUT_368E 16'h3636
`define CUBE_LUT_368F 16'h3637
`define CUBE_LUT_3690 16'h3638
`define CUBE_LUT_3691 16'h3639
`define CUBE_LUT_3692 16'h3639
`define CUBE_LUT_3693 16'h363A
`define CUBE_LUT_3694 16'h363B
`define CUBE_LUT_3695 16'h363C
`define CUBE_LUT_3696 16'h363D
`define CUBE_LUT_3697 16'h363E
`define CUBE_LUT_3698 16'h363F
`define CUBE_LUT_3699 16'h363F
`define CUBE_LUT_369A 16'h3640
`define CUBE_LUT_369B 16'h3641
`define CUBE_LUT_369C 16'h3642
`define CUBE_LUT_369D 16'h3643
`define CUBE_LUT_369E 16'h3644
`define CUBE_LUT_369F 16'h3644
`define CUBE_LUT_36A0 16'h3645
`define CUBE_LUT_36A1 16'h3646
`define CUBE_LUT_36A2 16'h3647
`define CUBE_LUT_36A3 16'h3648
`define CUBE_LUT_36A4 16'h3649
`define CUBE_LUT_36A5 16'h364A
`define CUBE_LUT_36A6 16'h364A
`define CUBE_LUT_36A7 16'h364B
`define CUBE_LUT_36A8 16'h364C
`define CUBE_LUT_36A9 16'h364D
`define CUBE_LUT_36AA 16'h364E
`define CUBE_LUT_36AB 16'h364F
`define CUBE_LUT_36AC 16'h364F
`define CUBE_LUT_36AD 16'h3650
`define CUBE_LUT_36AE 16'h3651
`define CUBE_LUT_36AF 16'h3652
`define CUBE_LUT_36B0 16'h3653
`define CUBE_LUT_36B1 16'h3654
`define CUBE_LUT_36B2 16'h3654
`define CUBE_LUT_36B3 16'h3655
`define CUBE_LUT_36B4 16'h3656
`define CUBE_LUT_36B5 16'h3657
`define CUBE_LUT_36B6 16'h3658
`define CUBE_LUT_36B7 16'h3659
`define CUBE_LUT_36B8 16'h365A
`define CUBE_LUT_36B9 16'h365A
`define CUBE_LUT_36BA 16'h365B
`define CUBE_LUT_36BB 16'h365C
`define CUBE_LUT_36BC 16'h365D
`define CUBE_LUT_36BD 16'h365E
`define CUBE_LUT_36BE 16'h365F
`define CUBE_LUT_36BF 16'h365F
`define CUBE_LUT_36C0 16'h3660
`define CUBE_LUT_36C1 16'h3661
`define CUBE_LUT_36C2 16'h3662
`define CUBE_LUT_36C3 16'h3663
`define CUBE_LUT_36C4 16'h3664
`define CUBE_LUT_36C5 16'h3664
`define CUBE_LUT_36C6 16'h3665
`define CUBE_LUT_36C7 16'h3666
`define CUBE_LUT_36C8 16'h3667
`define CUBE_LUT_36C9 16'h3668
`define CUBE_LUT_36CA 16'h3669
`define CUBE_LUT_36CB 16'h366A
`define CUBE_LUT_36CC 16'h366A
`define CUBE_LUT_36CD 16'h366B
`define CUBE_LUT_36CE 16'h366C
`define CUBE_LUT_36CF 16'h366D
`define CUBE_LUT_36D0 16'h366E
`define CUBE_LUT_36D1 16'h366F
`define CUBE_LUT_36D2 16'h366F
`define CUBE_LUT_36D3 16'h3670
`define CUBE_LUT_36D4 16'h3671
`define CUBE_LUT_36D5 16'h3672
`define CUBE_LUT_36D6 16'h3673
`define CUBE_LUT_36D7 16'h3674
`define CUBE_LUT_36D8 16'h3674
`define CUBE_LUT_36D9 16'h3675
`define CUBE_LUT_36DA 16'h3676
`define CUBE_LUT_36DB 16'h3677
`define CUBE_LUT_36DC 16'h3678
`define CUBE_LUT_36DD 16'h3679
`define CUBE_LUT_36DE 16'h3679
`define CUBE_LUT_36DF 16'h367A
`define CUBE_LUT_36E0 16'h367B
`define CUBE_LUT_36E1 16'h367C
`define CUBE_LUT_36E2 16'h367D
`define CUBE_LUT_36E3 16'h367E
`define CUBE_LUT_36E4 16'h367E
`define CUBE_LUT_36E5 16'h367F
`define CUBE_LUT_36E6 16'h3680
`define CUBE_LUT_36E7 16'h3681
`define CUBE_LUT_36E8 16'h3682
`define CUBE_LUT_36E9 16'h3683
`define CUBE_LUT_36EA 16'h3683
`define CUBE_LUT_36EB 16'h3684
`define CUBE_LUT_36EC 16'h3685
`define CUBE_LUT_36ED 16'h3686
`define CUBE_LUT_36EE 16'h3687
`define CUBE_LUT_36EF 16'h3688
`define CUBE_LUT_36F0 16'h3688
`define CUBE_LUT_36F1 16'h3689
`define CUBE_LUT_36F2 16'h368A
`define CUBE_LUT_36F3 16'h368B
`define CUBE_LUT_36F4 16'h368C
`define CUBE_LUT_36F5 16'h368D
`define CUBE_LUT_36F6 16'h368D
`define CUBE_LUT_36F7 16'h368E
`define CUBE_LUT_36F8 16'h368F
`define CUBE_LUT_36F9 16'h3690
`define CUBE_LUT_36FA 16'h3691
`define CUBE_LUT_36FB 16'h3692
`define CUBE_LUT_36FC 16'h3692
`define CUBE_LUT_36FD 16'h3693
`define CUBE_LUT_36FE 16'h3694
`define CUBE_LUT_36FF 16'h3695
`define CUBE_LUT_3700 16'h3696
`define CUBE_LUT_3701 16'h3697
`define CUBE_LUT_3702 16'h3697
`define CUBE_LUT_3703 16'h3698
`define CUBE_LUT_3704 16'h3699
`define CUBE_LUT_3705 16'h369A
`define CUBE_LUT_3706 16'h369B
`define CUBE_LUT_3707 16'h369C
`define CUBE_LUT_3708 16'h369C
`define CUBE_LUT_3709 16'h369D
`define CUBE_LUT_370A 16'h369E
`define CUBE_LUT_370B 16'h369F
`define CUBE_LUT_370C 16'h36A0
`define CUBE_LUT_370D 16'h36A1
`define CUBE_LUT_370E 16'h36A1
`define CUBE_LUT_370F 16'h36A2
`define CUBE_LUT_3710 16'h36A3
`define CUBE_LUT_3711 16'h36A4
`define CUBE_LUT_3712 16'h36A5
`define CUBE_LUT_3713 16'h36A6
`define CUBE_LUT_3714 16'h36A6
`define CUBE_LUT_3715 16'h36A7
`define CUBE_LUT_3716 16'h36A8
`define CUBE_LUT_3717 16'h36A9
`define CUBE_LUT_3718 16'h36AA
`define CUBE_LUT_3719 16'h36AB
`define CUBE_LUT_371A 16'h36AB
`define CUBE_LUT_371B 16'h36AC
`define CUBE_LUT_371C 16'h36AD
`define CUBE_LUT_371D 16'h36AE
`define CUBE_LUT_371E 16'h36AF
`define CUBE_LUT_371F 16'h36AF
`define CUBE_LUT_3720 16'h36B0
`define CUBE_LUT_3721 16'h36B1
`define CUBE_LUT_3722 16'h36B2
`define CUBE_LUT_3723 16'h36B3
`define CUBE_LUT_3724 16'h36B4
`define CUBE_LUT_3725 16'h36B4
`define CUBE_LUT_3726 16'h36B5
`define CUBE_LUT_3727 16'h36B6
`define CUBE_LUT_3728 16'h36B7
`define CUBE_LUT_3729 16'h36B8
`define CUBE_LUT_372A 16'h36B9
`define CUBE_LUT_372B 16'h36B9
`define CUBE_LUT_372C 16'h36BA
`define CUBE_LUT_372D 16'h36BB
`define CUBE_LUT_372E 16'h36BC
`define CUBE_LUT_372F 16'h36BD
`define CUBE_LUT_3730 16'h36BD
`define CUBE_LUT_3731 16'h36BE
`define CUBE_LUT_3732 16'h36BF
`define CUBE_LUT_3733 16'h36C0
`define CUBE_LUT_3734 16'h36C1
`define CUBE_LUT_3735 16'h36C2
`define CUBE_LUT_3736 16'h36C2
`define CUBE_LUT_3737 16'h36C3
`define CUBE_LUT_3738 16'h36C4
`define CUBE_LUT_3739 16'h36C5
`define CUBE_LUT_373A 16'h36C6
`define CUBE_LUT_373B 16'h36C7
`define CUBE_LUT_373C 16'h36C7
`define CUBE_LUT_373D 16'h36C8
`define CUBE_LUT_373E 16'h36C9
`define CUBE_LUT_373F 16'h36CA
`define CUBE_LUT_3740 16'h36CB
`define CUBE_LUT_3741 16'h36CB
`define CUBE_LUT_3742 16'h36CC
`define CUBE_LUT_3743 16'h36CD
`define CUBE_LUT_3744 16'h36CE
`define CUBE_LUT_3745 16'h36CF
`define CUBE_LUT_3746 16'h36D0
`define CUBE_LUT_3747 16'h36D0
`define CUBE_LUT_3748 16'h36D1
`define CUBE_LUT_3749 16'h36D2
`define CUBE_LUT_374A 16'h36D3
`define CUBE_LUT_374B 16'h36D4
`define CUBE_LUT_374C 16'h36D4
`define CUBE_LUT_374D 16'h36D5
`define CUBE_LUT_374E 16'h36D6
`define CUBE_LUT_374F 16'h36D7
`define CUBE_LUT_3750 16'h36D8
`define CUBE_LUT_3751 16'h36D9
`define CUBE_LUT_3752 16'h36D9
`define CUBE_LUT_3753 16'h36DA
`define CUBE_LUT_3754 16'h36DB
`define CUBE_LUT_3755 16'h36DC
`define CUBE_LUT_3756 16'h36DD
`define CUBE_LUT_3757 16'h36DD
`define CUBE_LUT_3758 16'h36DE
`define CUBE_LUT_3759 16'h36DF
`define CUBE_LUT_375A 16'h36E0
`define CUBE_LUT_375B 16'h36E1
`define CUBE_LUT_375C 16'h36E1
`define CUBE_LUT_375D 16'h36E2
`define CUBE_LUT_375E 16'h36E3
`define CUBE_LUT_375F 16'h36E4
`define CUBE_LUT_3760 16'h36E5
`define CUBE_LUT_3761 16'h36E6
`define CUBE_LUT_3762 16'h36E6
`define CUBE_LUT_3763 16'h36E7
`define CUBE_LUT_3764 16'h36E8
`define CUBE_LUT_3765 16'h36E9
`define CUBE_LUT_3766 16'h36EA
`define CUBE_LUT_3767 16'h36EA
`define CUBE_LUT_3768 16'h36EB
`define CUBE_LUT_3769 16'h36EC
`define CUBE_LUT_376A 16'h36ED
`define CUBE_LUT_376B 16'h36EE
`define CUBE_LUT_376C 16'h36EF
`define CUBE_LUT_376D 16'h36EF
`define CUBE_LUT_376E 16'h36F0
`define CUBE_LUT_376F 16'h36F1
`define CUBE_LUT_3770 16'h36F2
`define CUBE_LUT_3771 16'h36F3
`define CUBE_LUT_3772 16'h36F3
`define CUBE_LUT_3773 16'h36F4
`define CUBE_LUT_3774 16'h36F5
`define CUBE_LUT_3775 16'h36F6
`define CUBE_LUT_3776 16'h36F7
`define CUBE_LUT_3777 16'h36F7
`define CUBE_LUT_3778 16'h36F8
`define CUBE_LUT_3779 16'h36F9
`define CUBE_LUT_377A 16'h36FA
`define CUBE_LUT_377B 16'h36FB
`define CUBE_LUT_377C 16'h36FB
`define CUBE_LUT_377D 16'h36FC
`define CUBE_LUT_377E 16'h36FD
`define CUBE_LUT_377F 16'h36FE
`define CUBE_LUT_3780 16'h36FF
`define CUBE_LUT_3781 16'h3700
`define CUBE_LUT_3782 16'h3700
`define CUBE_LUT_3783 16'h3701
`define CUBE_LUT_3784 16'h3702
`define CUBE_LUT_3785 16'h3703
`define CUBE_LUT_3786 16'h3704
`define CUBE_LUT_3787 16'h3704
`define CUBE_LUT_3788 16'h3705
`define CUBE_LUT_3789 16'h3706
`define CUBE_LUT_378A 16'h3707
`define CUBE_LUT_378B 16'h3708
`define CUBE_LUT_378C 16'h3708
`define CUBE_LUT_378D 16'h3709
`define CUBE_LUT_378E 16'h370A
`define CUBE_LUT_378F 16'h370B
`define CUBE_LUT_3790 16'h370C
`define CUBE_LUT_3791 16'h370C
`define CUBE_LUT_3792 16'h370D
`define CUBE_LUT_3793 16'h370E
`define CUBE_LUT_3794 16'h370F
`define CUBE_LUT_3795 16'h3710
`define CUBE_LUT_3796 16'h3710
`define CUBE_LUT_3797 16'h3711
`define CUBE_LUT_3798 16'h3712
`define CUBE_LUT_3799 16'h3713
`define CUBE_LUT_379A 16'h3714
`define CUBE_LUT_379B 16'h3715
`define CUBE_LUT_379C 16'h3715
`define CUBE_LUT_379D 16'h3716
`define CUBE_LUT_379E 16'h3717
`define CUBE_LUT_379F 16'h3718
`define CUBE_LUT_37A0 16'h3719
`define CUBE_LUT_37A1 16'h3719
`define CUBE_LUT_37A2 16'h371A
`define CUBE_LUT_37A3 16'h371B
`define CUBE_LUT_37A4 16'h371C
`define CUBE_LUT_37A5 16'h371D
`define CUBE_LUT_37A6 16'h371D
`define CUBE_LUT_37A7 16'h371E
`define CUBE_LUT_37A8 16'h371F
`define CUBE_LUT_37A9 16'h3720
`define CUBE_LUT_37AA 16'h3721
`define CUBE_LUT_37AB 16'h3721
`define CUBE_LUT_37AC 16'h3722
`define CUBE_LUT_37AD 16'h3723
`define CUBE_LUT_37AE 16'h3724
`define CUBE_LUT_37AF 16'h3725
`define CUBE_LUT_37B0 16'h3725
`define CUBE_LUT_37B1 16'h3726
`define CUBE_LUT_37B2 16'h3727
`define CUBE_LUT_37B3 16'h3728
`define CUBE_LUT_37B4 16'h3729
`define CUBE_LUT_37B5 16'h3729
`define CUBE_LUT_37B6 16'h372A
`define CUBE_LUT_37B7 16'h372B
`define CUBE_LUT_37B8 16'h372C
`define CUBE_LUT_37B9 16'h372D
`define CUBE_LUT_37BA 16'h372D
`define CUBE_LUT_37BB 16'h372E
`define CUBE_LUT_37BC 16'h372F
`define CUBE_LUT_37BD 16'h3730
`define CUBE_LUT_37BE 16'h3731
`define CUBE_LUT_37BF 16'h3731
`define CUBE_LUT_37C0 16'h3732
`define CUBE_LUT_37C1 16'h3733
`define CUBE_LUT_37C2 16'h3734
`define CUBE_LUT_37C3 16'h3735
`define CUBE_LUT_37C4 16'h3735
`define CUBE_LUT_37C5 16'h3736
`define CUBE_LUT_37C6 16'h3737
`define CUBE_LUT_37C7 16'h3738
`define CUBE_LUT_37C8 16'h3739
`define CUBE_LUT_37C9 16'h3739
`define CUBE_LUT_37CA 16'h373A
`define CUBE_LUT_37CB 16'h373B
`define CUBE_LUT_37CC 16'h373C
`define CUBE_LUT_37CD 16'h373C
`define CUBE_LUT_37CE 16'h373D
`define CUBE_LUT_37CF 16'h373E
`define CUBE_LUT_37D0 16'h373F
`define CUBE_LUT_37D1 16'h3740
`define CUBE_LUT_37D2 16'h3740
`define CUBE_LUT_37D3 16'h3741
`define CUBE_LUT_37D4 16'h3742
`define CUBE_LUT_37D5 16'h3743
`define CUBE_LUT_37D6 16'h3744
`define CUBE_LUT_37D7 16'h3744
`define CUBE_LUT_37D8 16'h3745
`define CUBE_LUT_37D9 16'h3746
`define CUBE_LUT_37DA 16'h3747
`define CUBE_LUT_37DB 16'h3748
`define CUBE_LUT_37DC 16'h3748
`define CUBE_LUT_37DD 16'h3749
`define CUBE_LUT_37DE 16'h374A
`define CUBE_LUT_37DF 16'h374B
`define CUBE_LUT_37E0 16'h374C
`define CUBE_LUT_37E1 16'h374C
`define CUBE_LUT_37E2 16'h374D
`define CUBE_LUT_37E3 16'h374E
`define CUBE_LUT_37E4 16'h374F
`define CUBE_LUT_37E5 16'h3750
`define CUBE_LUT_37E6 16'h3750
`define CUBE_LUT_37E7 16'h3751
`define CUBE_LUT_37E8 16'h3752
`define CUBE_LUT_37E9 16'h3753
`define CUBE_LUT_37EA 16'h3753
`define CUBE_LUT_37EB 16'h3754
`define CUBE_LUT_37EC 16'h3755
`define CUBE_LUT_37ED 16'h3756
`define CUBE_LUT_37EE 16'h3757
`define CUBE_LUT_37EF 16'h3757
`define CUBE_LUT_37F0 16'h3758
`define CUBE_LUT_37F1 16'h3759
`define CUBE_LUT_37F2 16'h375A
`define CUBE_LUT_37F3 16'h375B
`define CUBE_LUT_37F4 16'h375B
`define CUBE_LUT_37F5 16'h375C
`define CUBE_LUT_37F6 16'h375D
`define CUBE_LUT_37F7 16'h375E
`define CUBE_LUT_37F8 16'h375F
`define CUBE_LUT_37F9 16'h375F
`define CUBE_LUT_37FA 16'h3760
`define CUBE_LUT_37FB 16'h3761
`define CUBE_LUT_37FC 16'h3762
`define CUBE_LUT_37FD 16'h3762
`define CUBE_LUT_37FE 16'h3763
`define CUBE_LUT_37FF 16'h3764
`define CUBE_LUT_3800 16'h3765
`define CUBE_LUT_3801 16'h3766
`define CUBE_LUT_3802 16'h3768
`define CUBE_LUT_3803 16'h376A
`define CUBE_LUT_3804 16'h376B
`define CUBE_LUT_3805 16'h376D
`define CUBE_LUT_3806 16'h376E
`define CUBE_LUT_3807 16'h3770
`define CUBE_LUT_3808 16'h3771
`define CUBE_LUT_3809 16'h3773
`define CUBE_LUT_380A 16'h3775
`define CUBE_LUT_380B 16'h3776
`define CUBE_LUT_380C 16'h3778
`define CUBE_LUT_380D 16'h3779
`define CUBE_LUT_380E 16'h377B
`define CUBE_LUT_380F 16'h377C
`define CUBE_LUT_3810 16'h377E
`define CUBE_LUT_3811 16'h377F
`define CUBE_LUT_3812 16'h3781
`define CUBE_LUT_3813 16'h3783
`define CUBE_LUT_3814 16'h3784
`define CUBE_LUT_3815 16'h3786
`define CUBE_LUT_3816 16'h3787
`define CUBE_LUT_3817 16'h3789
`define CUBE_LUT_3818 16'h378A
`define CUBE_LUT_3819 16'h378C
`define CUBE_LUT_381A 16'h378D
`define CUBE_LUT_381B 16'h378F
`define CUBE_LUT_381C 16'h3791
`define CUBE_LUT_381D 16'h3792
`define CUBE_LUT_381E 16'h3794
`define CUBE_LUT_381F 16'h3795
`define CUBE_LUT_3820 16'h3797
`define CUBE_LUT_3821 16'h3798
`define CUBE_LUT_3822 16'h379A
`define CUBE_LUT_3823 16'h379B
`define CUBE_LUT_3824 16'h379D
`define CUBE_LUT_3825 16'h379F
`define CUBE_LUT_3826 16'h37A0
`define CUBE_LUT_3827 16'h37A2
`define CUBE_LUT_3828 16'h37A3
`define CUBE_LUT_3829 16'h37A5
`define CUBE_LUT_382A 16'h37A6
`define CUBE_LUT_382B 16'h37A8
`define CUBE_LUT_382C 16'h37A9
`define CUBE_LUT_382D 16'h37AB
`define CUBE_LUT_382E 16'h37AC
`define CUBE_LUT_382F 16'h37AE
`define CUBE_LUT_3830 16'h37B0
`define CUBE_LUT_3831 16'h37B1
`define CUBE_LUT_3832 16'h37B3
`define CUBE_LUT_3833 16'h37B4
`define CUBE_LUT_3834 16'h37B6
`define CUBE_LUT_3835 16'h37B7
`define CUBE_LUT_3836 16'h37B9
`define CUBE_LUT_3837 16'h37BA
`define CUBE_LUT_3838 16'h37BC
`define CUBE_LUT_3839 16'h37BD
`define CUBE_LUT_383A 16'h37BF
`define CUBE_LUT_383B 16'h37C0
`define CUBE_LUT_383C 16'h37C2
`define CUBE_LUT_383D 16'h37C3
`define CUBE_LUT_383E 16'h37C5
`define CUBE_LUT_383F 16'h37C7
`define CUBE_LUT_3840 16'h37C8
`define CUBE_LUT_3841 16'h37CA
`define CUBE_LUT_3842 16'h37CB
`define CUBE_LUT_3843 16'h37CD
`define CUBE_LUT_3844 16'h37CE
`define CUBE_LUT_3845 16'h37D0
`define CUBE_LUT_3846 16'h37D1
`define CUBE_LUT_3847 16'h37D3
`define CUBE_LUT_3848 16'h37D4
`define CUBE_LUT_3849 16'h37D6
`define CUBE_LUT_384A 16'h37D7
`define CUBE_LUT_384B 16'h37D9
`define CUBE_LUT_384C 16'h37DA
`define CUBE_LUT_384D 16'h37DC
`define CUBE_LUT_384E 16'h37DD
`define CUBE_LUT_384F 16'h37DF
`define CUBE_LUT_3850 16'h37E0
`define CUBE_LUT_3851 16'h37E2
`define CUBE_LUT_3852 16'h37E3
`define CUBE_LUT_3853 16'h37E5
`define CUBE_LUT_3854 16'h37E6
`define CUBE_LUT_3855 16'h37E8
`define CUBE_LUT_3856 16'h37E9
`define CUBE_LUT_3857 16'h37EB
`define CUBE_LUT_3858 16'h37EC
`define CUBE_LUT_3859 16'h37EE
`define CUBE_LUT_385A 16'h37EF
`define CUBE_LUT_385B 16'h37F1
`define CUBE_LUT_385C 16'h37F3
`define CUBE_LUT_385D 16'h37F4
`define CUBE_LUT_385E 16'h37F6
`define CUBE_LUT_385F 16'h37F7
`define CUBE_LUT_3860 16'h37F9
`define CUBE_LUT_3861 16'h37FA
`define CUBE_LUT_3862 16'h37FC
`define CUBE_LUT_3863 16'h37FD
`define CUBE_LUT_3864 16'h37FF
`define CUBE_LUT_3865 16'h3800
`define CUBE_LUT_3866 16'h3801
`define CUBE_LUT_3867 16'h3802
`define CUBE_LUT_3868 16'h3802
`define CUBE_LUT_3869 16'h3803
`define CUBE_LUT_386A 16'h3804
`define CUBE_LUT_386B 16'h3805
`define CUBE_LUT_386C 16'h3805
`define CUBE_LUT_386D 16'h3806
`define CUBE_LUT_386E 16'h3807
`define CUBE_LUT_386F 16'h3807
`define CUBE_LUT_3870 16'h3808
`define CUBE_LUT_3871 16'h3809
`define CUBE_LUT_3872 16'h380A
`define CUBE_LUT_3873 16'h380A
`define CUBE_LUT_3874 16'h380B
`define CUBE_LUT_3875 16'h380C
`define CUBE_LUT_3876 16'h380D
`define CUBE_LUT_3877 16'h380D
`define CUBE_LUT_3878 16'h380E
`define CUBE_LUT_3879 16'h380F
`define CUBE_LUT_387A 16'h3810
`define CUBE_LUT_387B 16'h3810
`define CUBE_LUT_387C 16'h3811
`define CUBE_LUT_387D 16'h3812
`define CUBE_LUT_387E 16'h3813
`define CUBE_LUT_387F 16'h3813
`define CUBE_LUT_3880 16'h3814
`define CUBE_LUT_3881 16'h3815
`define CUBE_LUT_3882 16'h3816
`define CUBE_LUT_3883 16'h3816
`define CUBE_LUT_3884 16'h3817
`define CUBE_LUT_3885 16'h3818
`define CUBE_LUT_3886 16'h3819
`define CUBE_LUT_3887 16'h3819
`define CUBE_LUT_3888 16'h381A
`define CUBE_LUT_3889 16'h381B
`define CUBE_LUT_388A 16'h381C
`define CUBE_LUT_388B 16'h381C
`define CUBE_LUT_388C 16'h381D
`define CUBE_LUT_388D 16'h381E
`define CUBE_LUT_388E 16'h381E
`define CUBE_LUT_388F 16'h381F
`define CUBE_LUT_3890 16'h3820
`define CUBE_LUT_3891 16'h3821
`define CUBE_LUT_3892 16'h3821
`define CUBE_LUT_3893 16'h3822
`define CUBE_LUT_3894 16'h3823
`define CUBE_LUT_3895 16'h3824
`define CUBE_LUT_3896 16'h3824
`define CUBE_LUT_3897 16'h3825
`define CUBE_LUT_3898 16'h3826
`define CUBE_LUT_3899 16'h3827
`define CUBE_LUT_389A 16'h3827
`define CUBE_LUT_389B 16'h3828
`define CUBE_LUT_389C 16'h3829
`define CUBE_LUT_389D 16'h3829
`define CUBE_LUT_389E 16'h382A
`define CUBE_LUT_389F 16'h382B
`define CUBE_LUT_38A0 16'h382C
`define CUBE_LUT_38A1 16'h382C
`define CUBE_LUT_38A2 16'h382D
`define CUBE_LUT_38A3 16'h382E
`define CUBE_LUT_38A4 16'h382F
`define CUBE_LUT_38A5 16'h382F
`define CUBE_LUT_38A6 16'h3830
`define CUBE_LUT_38A7 16'h3831
`define CUBE_LUT_38A8 16'h3831
`define CUBE_LUT_38A9 16'h3832
`define CUBE_LUT_38AA 16'h3833
`define CUBE_LUT_38AB 16'h3834
`define CUBE_LUT_38AC 16'h3834
`define CUBE_LUT_38AD 16'h3835
`define CUBE_LUT_38AE 16'h3836
`define CUBE_LUT_38AF 16'h3837
`define CUBE_LUT_38B0 16'h3837
`define CUBE_LUT_38B1 16'h3838
`define CUBE_LUT_38B2 16'h3839
`define CUBE_LUT_38B3 16'h3839
`define CUBE_LUT_38B4 16'h383A
`define CUBE_LUT_38B5 16'h383B
`define CUBE_LUT_38B6 16'h383C
`define CUBE_LUT_38B7 16'h383C
`define CUBE_LUT_38B8 16'h383D
`define CUBE_LUT_38B9 16'h383E
`define CUBE_LUT_38BA 16'h383E
`define CUBE_LUT_38BB 16'h383F
`define CUBE_LUT_38BC 16'h3840
`define CUBE_LUT_38BD 16'h3841
`define CUBE_LUT_38BE 16'h3841
`define CUBE_LUT_38BF 16'h3842
`define CUBE_LUT_38C0 16'h3843
`define CUBE_LUT_38C1 16'h3843
`define CUBE_LUT_38C2 16'h3844
`define CUBE_LUT_38C3 16'h3845
`define CUBE_LUT_38C4 16'h3846
`define CUBE_LUT_38C5 16'h3846
`define CUBE_LUT_38C6 16'h3847
`define CUBE_LUT_38C7 16'h3848
`define CUBE_LUT_38C8 16'h3848
`define CUBE_LUT_38C9 16'h3849
`define CUBE_LUT_38CA 16'h384A
`define CUBE_LUT_38CB 16'h384B
`define CUBE_LUT_38CC 16'h384B
`define CUBE_LUT_38CD 16'h384C
`define CUBE_LUT_38CE 16'h384D
`define CUBE_LUT_38CF 16'h384D
`define CUBE_LUT_38D0 16'h384E
`define CUBE_LUT_38D1 16'h384F
`define CUBE_LUT_38D2 16'h3850
`define CUBE_LUT_38D3 16'h3850
`define CUBE_LUT_38D4 16'h3851
`define CUBE_LUT_38D5 16'h3852
`define CUBE_LUT_38D6 16'h3852
`define CUBE_LUT_38D7 16'h3853
`define CUBE_LUT_38D8 16'h3854
`define CUBE_LUT_38D9 16'h3855
`define CUBE_LUT_38DA 16'h3855
`define CUBE_LUT_38DB 16'h3856
`define CUBE_LUT_38DC 16'h3857
`define CUBE_LUT_38DD 16'h3857
`define CUBE_LUT_38DE 16'h3858
`define CUBE_LUT_38DF 16'h3859
`define CUBE_LUT_38E0 16'h3859
`define CUBE_LUT_38E1 16'h385A
`define CUBE_LUT_38E2 16'h385B
`define CUBE_LUT_38E3 16'h385C
`define CUBE_LUT_38E4 16'h385C
`define CUBE_LUT_38E5 16'h385D
`define CUBE_LUT_38E6 16'h385E
`define CUBE_LUT_38E7 16'h385E
`define CUBE_LUT_38E8 16'h385F
`define CUBE_LUT_38E9 16'h3860
`define CUBE_LUT_38EA 16'h3860
`define CUBE_LUT_38EB 16'h3861
`define CUBE_LUT_38EC 16'h3862
`define CUBE_LUT_38ED 16'h3863
`define CUBE_LUT_38EE 16'h3863
`define CUBE_LUT_38EF 16'h3864
`define CUBE_LUT_38F0 16'h3865
`define CUBE_LUT_38F1 16'h3865
`define CUBE_LUT_38F2 16'h3866
`define CUBE_LUT_38F3 16'h3867
`define CUBE_LUT_38F4 16'h3867
`define CUBE_LUT_38F5 16'h3868
`define CUBE_LUT_38F6 16'h3869
`define CUBE_LUT_38F7 16'h386A
`define CUBE_LUT_38F8 16'h386A
`define CUBE_LUT_38F9 16'h386B
`define CUBE_LUT_38FA 16'h386C
`define CUBE_LUT_38FB 16'h386C
`define CUBE_LUT_38FC 16'h386D
`define CUBE_LUT_38FD 16'h386E
`define CUBE_LUT_38FE 16'h386E
`define CUBE_LUT_38FF 16'h386F
`define CUBE_LUT_3900 16'h3870
`define CUBE_LUT_3901 16'h3871
`define CUBE_LUT_3902 16'h3871
`define CUBE_LUT_3903 16'h3872
`define CUBE_LUT_3904 16'h3873
`define CUBE_LUT_3905 16'h3873
`define CUBE_LUT_3906 16'h3874
`define CUBE_LUT_3907 16'h3875
`define CUBE_LUT_3908 16'h3875
`define CUBE_LUT_3909 16'h3876
`define CUBE_LUT_390A 16'h3877
`define CUBE_LUT_390B 16'h3877
`define CUBE_LUT_390C 16'h3878
`define CUBE_LUT_390D 16'h3879
`define CUBE_LUT_390E 16'h3879
`define CUBE_LUT_390F 16'h387A
`define CUBE_LUT_3910 16'h387B
`define CUBE_LUT_3911 16'h387C
`define CUBE_LUT_3912 16'h387C
`define CUBE_LUT_3913 16'h387D
`define CUBE_LUT_3914 16'h387E
`define CUBE_LUT_3915 16'h387E
`define CUBE_LUT_3916 16'h387F
`define CUBE_LUT_3917 16'h3880
`define CUBE_LUT_3918 16'h3880
`define CUBE_LUT_3919 16'h3881
`define CUBE_LUT_391A 16'h3882
`define CUBE_LUT_391B 16'h3882
`define CUBE_LUT_391C 16'h3883
`define CUBE_LUT_391D 16'h3884
`define CUBE_LUT_391E 16'h3884
`define CUBE_LUT_391F 16'h3885
`define CUBE_LUT_3920 16'h3886
`define CUBE_LUT_3921 16'h3886
`define CUBE_LUT_3922 16'h3887
`define CUBE_LUT_3923 16'h3888
`define CUBE_LUT_3924 16'h3889
`define CUBE_LUT_3925 16'h3889
`define CUBE_LUT_3926 16'h388A
`define CUBE_LUT_3927 16'h388B
`define CUBE_LUT_3928 16'h388B
`define CUBE_LUT_3929 16'h388C
`define CUBE_LUT_392A 16'h388D
`define CUBE_LUT_392B 16'h388D
`define CUBE_LUT_392C 16'h388E
`define CUBE_LUT_392D 16'h388F
`define CUBE_LUT_392E 16'h388F
`define CUBE_LUT_392F 16'h3890
`define CUBE_LUT_3930 16'h3891
`define CUBE_LUT_3931 16'h3891
`define CUBE_LUT_3932 16'h3892
`define CUBE_LUT_3933 16'h3893
`define CUBE_LUT_3934 16'h3893
`define CUBE_LUT_3935 16'h3894
`define CUBE_LUT_3936 16'h3895
`define CUBE_LUT_3937 16'h3895
`define CUBE_LUT_3938 16'h3896
`define CUBE_LUT_3939 16'h3897
`define CUBE_LUT_393A 16'h3897
`define CUBE_LUT_393B 16'h3898
`define CUBE_LUT_393C 16'h3899
`define CUBE_LUT_393D 16'h3899
`define CUBE_LUT_393E 16'h389A
`define CUBE_LUT_393F 16'h389B
`define CUBE_LUT_3940 16'h389B
`define CUBE_LUT_3941 16'h389C
`define CUBE_LUT_3942 16'h389D
`define CUBE_LUT_3943 16'h389D
`define CUBE_LUT_3944 16'h389E
`define CUBE_LUT_3945 16'h389F
`define CUBE_LUT_3946 16'h389F
`define CUBE_LUT_3947 16'h38A0
`define CUBE_LUT_3948 16'h38A1
`define CUBE_LUT_3949 16'h38A1
`define CUBE_LUT_394A 16'h38A2
`define CUBE_LUT_394B 16'h38A3
`define CUBE_LUT_394C 16'h38A3
`define CUBE_LUT_394D 16'h38A4
`define CUBE_LUT_394E 16'h38A5
`define CUBE_LUT_394F 16'h38A5
`define CUBE_LUT_3950 16'h38A6
`define CUBE_LUT_3951 16'h38A7
`define CUBE_LUT_3952 16'h38A7
`define CUBE_LUT_3953 16'h38A8
`define CUBE_LUT_3954 16'h38A9
`define CUBE_LUT_3955 16'h38A9
`define CUBE_LUT_3956 16'h38AA
`define CUBE_LUT_3957 16'h38AB
`define CUBE_LUT_3958 16'h38AB
`define CUBE_LUT_3959 16'h38AC
`define CUBE_LUT_395A 16'h38AD
`define CUBE_LUT_395B 16'h38AD
`define CUBE_LUT_395C 16'h38AE
`define CUBE_LUT_395D 16'h38AF
`define CUBE_LUT_395E 16'h38AF
`define CUBE_LUT_395F 16'h38B0
`define CUBE_LUT_3960 16'h38B1
`define CUBE_LUT_3961 16'h38B1
`define CUBE_LUT_3962 16'h38B2
`define CUBE_LUT_3963 16'h38B3
`define CUBE_LUT_3964 16'h38B3
`define CUBE_LUT_3965 16'h38B4
`define CUBE_LUT_3966 16'h38B4
`define CUBE_LUT_3967 16'h38B5
`define CUBE_LUT_3968 16'h38B6
`define CUBE_LUT_3969 16'h38B6
`define CUBE_LUT_396A 16'h38B7
`define CUBE_LUT_396B 16'h38B8
`define CUBE_LUT_396C 16'h38B8
`define CUBE_LUT_396D 16'h38B9
`define CUBE_LUT_396E 16'h38BA
`define CUBE_LUT_396F 16'h38BA
`define CUBE_LUT_3970 16'h38BB
`define CUBE_LUT_3971 16'h38BC
`define CUBE_LUT_3972 16'h38BC
`define CUBE_LUT_3973 16'h38BD
`define CUBE_LUT_3974 16'h38BE
`define CUBE_LUT_3975 16'h38BE
`define CUBE_LUT_3976 16'h38BF
`define CUBE_LUT_3977 16'h38C0
`define CUBE_LUT_3978 16'h38C0
`define CUBE_LUT_3979 16'h38C1
`define CUBE_LUT_397A 16'h38C2
`define CUBE_LUT_397B 16'h38C2
`define CUBE_LUT_397C 16'h38C3
`define CUBE_LUT_397D 16'h38C3
`define CUBE_LUT_397E 16'h38C4
`define CUBE_LUT_397F 16'h38C5
`define CUBE_LUT_3980 16'h38C5
`define CUBE_LUT_3981 16'h38C6
`define CUBE_LUT_3982 16'h38C7
`define CUBE_LUT_3983 16'h38C7
`define CUBE_LUT_3984 16'h38C8
`define CUBE_LUT_3985 16'h38C9
`define CUBE_LUT_3986 16'h38C9
`define CUBE_LUT_3987 16'h38CA
`define CUBE_LUT_3988 16'h38CB
`define CUBE_LUT_3989 16'h38CB
`define CUBE_LUT_398A 16'h38CC
`define CUBE_LUT_398B 16'h38CC
`define CUBE_LUT_398C 16'h38CD
`define CUBE_LUT_398D 16'h38CE
`define CUBE_LUT_398E 16'h38CE
`define CUBE_LUT_398F 16'h38CF
`define CUBE_LUT_3990 16'h38D0
`define CUBE_LUT_3991 16'h38D0
`define CUBE_LUT_3992 16'h38D1
`define CUBE_LUT_3993 16'h38D2
`define CUBE_LUT_3994 16'h38D2
`define CUBE_LUT_3995 16'h38D3
`define CUBE_LUT_3996 16'h38D3
`define CUBE_LUT_3997 16'h38D4
`define CUBE_LUT_3998 16'h38D5
`define CUBE_LUT_3999 16'h38D5
`define CUBE_LUT_399A 16'h38D6
`define CUBE_LUT_399B 16'h38D7
`define CUBE_LUT_399C 16'h38D7
`define CUBE_LUT_399D 16'h38D8
`define CUBE_LUT_399E 16'h38D9
`define CUBE_LUT_399F 16'h38D9
`define CUBE_LUT_39A0 16'h38DA
`define CUBE_LUT_39A1 16'h38DA
`define CUBE_LUT_39A2 16'h38DB
`define CUBE_LUT_39A3 16'h38DC
`define CUBE_LUT_39A4 16'h38DC
`define CUBE_LUT_39A5 16'h38DD
`define CUBE_LUT_39A6 16'h38DE
`define CUBE_LUT_39A7 16'h38DE
`define CUBE_LUT_39A8 16'h38DF
`define CUBE_LUT_39A9 16'h38DF
`define CUBE_LUT_39AA 16'h38E0
`define CUBE_LUT_39AB 16'h38E1
`define CUBE_LUT_39AC 16'h38E1
`define CUBE_LUT_39AD 16'h38E2
`define CUBE_LUT_39AE 16'h38E3
`define CUBE_LUT_39AF 16'h38E3
`define CUBE_LUT_39B0 16'h38E4
`define CUBE_LUT_39B1 16'h38E4
`define CUBE_LUT_39B2 16'h38E5
`define CUBE_LUT_39B3 16'h38E6
`define CUBE_LUT_39B4 16'h38E6
`define CUBE_LUT_39B5 16'h38E7
`define CUBE_LUT_39B6 16'h38E8
`define CUBE_LUT_39B7 16'h38E8
`define CUBE_LUT_39B8 16'h38E9
`define CUBE_LUT_39B9 16'h38E9
`define CUBE_LUT_39BA 16'h38EA
`define CUBE_LUT_39BB 16'h38EB
`define CUBE_LUT_39BC 16'h38EB
`define CUBE_LUT_39BD 16'h38EC
`define CUBE_LUT_39BE 16'h38ED
`define CUBE_LUT_39BF 16'h38ED
`define CUBE_LUT_39C0 16'h38EE
`define CUBE_LUT_39C1 16'h38EE
`define CUBE_LUT_39C2 16'h38EF
`define CUBE_LUT_39C3 16'h38F0
`define CUBE_LUT_39C4 16'h38F0
`define CUBE_LUT_39C5 16'h38F1
`define CUBE_LUT_39C6 16'h38F2
`define CUBE_LUT_39C7 16'h38F2
`define CUBE_LUT_39C8 16'h38F3
`define CUBE_LUT_39C9 16'h38F3
`define CUBE_LUT_39CA 16'h38F4
`define CUBE_LUT_39CB 16'h38F5
`define CUBE_LUT_39CC 16'h38F5
`define CUBE_LUT_39CD 16'h38F6
`define CUBE_LUT_39CE 16'h38F6
`define CUBE_LUT_39CF 16'h38F7
`define CUBE_LUT_39D0 16'h38F8
`define CUBE_LUT_39D1 16'h38F8
`define CUBE_LUT_39D2 16'h38F9
`define CUBE_LUT_39D3 16'h38FA
`define CUBE_LUT_39D4 16'h38FA
`define CUBE_LUT_39D5 16'h38FB
`define CUBE_LUT_39D6 16'h38FB
`define CUBE_LUT_39D7 16'h38FC
`define CUBE_LUT_39D8 16'h38FD
`define CUBE_LUT_39D9 16'h38FD
`define CUBE_LUT_39DA 16'h38FE
`define CUBE_LUT_39DB 16'h38FE
`define CUBE_LUT_39DC 16'h38FF
`define CUBE_LUT_39DD 16'h3900
`define CUBE_LUT_39DE 16'h3900
`define CUBE_LUT_39DF 16'h3901
`define CUBE_LUT_39E0 16'h3902
`define CUBE_LUT_39E1 16'h3902
`define CUBE_LUT_39E2 16'h3903
`define CUBE_LUT_39E3 16'h3903
`define CUBE_LUT_39E4 16'h3904
`define CUBE_LUT_39E5 16'h3905
`define CUBE_LUT_39E6 16'h3905
`define CUBE_LUT_39E7 16'h3906
`define CUBE_LUT_39E8 16'h3906
`define CUBE_LUT_39E9 16'h3907
`define CUBE_LUT_39EA 16'h3908
`define CUBE_LUT_39EB 16'h3908
`define CUBE_LUT_39EC 16'h3909
`define CUBE_LUT_39ED 16'h3909
`define CUBE_LUT_39EE 16'h390A
`define CUBE_LUT_39EF 16'h390B
`define CUBE_LUT_39F0 16'h390B
`define CUBE_LUT_39F1 16'h390C
`define CUBE_LUT_39F2 16'h390C
`define CUBE_LUT_39F3 16'h390D
`define CUBE_LUT_39F4 16'h390E
`define CUBE_LUT_39F5 16'h390E
`define CUBE_LUT_39F6 16'h390F
`define CUBE_LUT_39F7 16'h390F
`define CUBE_LUT_39F8 16'h3910
`define CUBE_LUT_39F9 16'h3911
`define CUBE_LUT_39FA 16'h3911
`define CUBE_LUT_39FB 16'h3912
`define CUBE_LUT_39FC 16'h3912
`define CUBE_LUT_39FD 16'h3913
`define CUBE_LUT_39FE 16'h3914
`define CUBE_LUT_39FF 16'h3914
`define CUBE_LUT_3A00 16'h3915
`define CUBE_LUT_3A01 16'h3915
`define CUBE_LUT_3A02 16'h3916
`define CUBE_LUT_3A03 16'h3917
`define CUBE_LUT_3A04 16'h3917
`define CUBE_LUT_3A05 16'h3918
`define CUBE_LUT_3A06 16'h3918
`define CUBE_LUT_3A07 16'h3919
`define CUBE_LUT_3A08 16'h391A
`define CUBE_LUT_3A09 16'h391A
`define CUBE_LUT_3A0A 16'h391B
`define CUBE_LUT_3A0B 16'h391B
`define CUBE_LUT_3A0C 16'h391C
`define CUBE_LUT_3A0D 16'h391D
`define CUBE_LUT_3A0E 16'h391D
`define CUBE_LUT_3A0F 16'h391E
`define CUBE_LUT_3A10 16'h391E
`define CUBE_LUT_3A11 16'h391F
`define CUBE_LUT_3A12 16'h391F
`define CUBE_LUT_3A13 16'h3920
`define CUBE_LUT_3A14 16'h3921
`define CUBE_LUT_3A15 16'h3921
`define CUBE_LUT_3A16 16'h3922
`define CUBE_LUT_3A17 16'h3922
`define CUBE_LUT_3A18 16'h3923
`define CUBE_LUT_3A19 16'h3924
`define CUBE_LUT_3A1A 16'h3924
`define CUBE_LUT_3A1B 16'h3925
`define CUBE_LUT_3A1C 16'h3925
`define CUBE_LUT_3A1D 16'h3926
`define CUBE_LUT_3A1E 16'h3927
`define CUBE_LUT_3A1F 16'h3927
`define CUBE_LUT_3A20 16'h3928
`define CUBE_LUT_3A21 16'h3928
`define CUBE_LUT_3A22 16'h3929
`define CUBE_LUT_3A23 16'h3929
`define CUBE_LUT_3A24 16'h392A
`define CUBE_LUT_3A25 16'h392B
`define CUBE_LUT_3A26 16'h392B
`define CUBE_LUT_3A27 16'h392C
`define CUBE_LUT_3A28 16'h392C
`define CUBE_LUT_3A29 16'h392D
`define CUBE_LUT_3A2A 16'h392E
`define CUBE_LUT_3A2B 16'h392E
`define CUBE_LUT_3A2C 16'h392F
`define CUBE_LUT_3A2D 16'h392F
`define CUBE_LUT_3A2E 16'h3930
`define CUBE_LUT_3A2F 16'h3930
`define CUBE_LUT_3A30 16'h3931
`define CUBE_LUT_3A31 16'h3932
`define CUBE_LUT_3A32 16'h3932
`define CUBE_LUT_3A33 16'h3933
`define CUBE_LUT_3A34 16'h3933
`define CUBE_LUT_3A35 16'h3934
`define CUBE_LUT_3A36 16'h3934
`define CUBE_LUT_3A37 16'h3935
`define CUBE_LUT_3A38 16'h3936
`define CUBE_LUT_3A39 16'h3936
`define CUBE_LUT_3A3A 16'h3937
`define CUBE_LUT_3A3B 16'h3937
`define CUBE_LUT_3A3C 16'h3938
`define CUBE_LUT_3A3D 16'h3938
`define CUBE_LUT_3A3E 16'h3939
`define CUBE_LUT_3A3F 16'h393A
`define CUBE_LUT_3A40 16'h393A
`define CUBE_LUT_3A41 16'h393B
`define CUBE_LUT_3A42 16'h393B
`define CUBE_LUT_3A43 16'h393C
`define CUBE_LUT_3A44 16'h393D
`define CUBE_LUT_3A45 16'h393D
`define CUBE_LUT_3A46 16'h393E
`define CUBE_LUT_3A47 16'h393E
`define CUBE_LUT_3A48 16'h393F
`define CUBE_LUT_3A49 16'h393F
`define CUBE_LUT_3A4A 16'h3940
`define CUBE_LUT_3A4B 16'h3940
`define CUBE_LUT_3A4C 16'h3941
`define CUBE_LUT_3A4D 16'h3942
`define CUBE_LUT_3A4E 16'h3942
`define CUBE_LUT_3A4F 16'h3943
`define CUBE_LUT_3A50 16'h3943
`define CUBE_LUT_3A51 16'h3944
`define CUBE_LUT_3A52 16'h3944
`define CUBE_LUT_3A53 16'h3945
`define CUBE_LUT_3A54 16'h3946
`define CUBE_LUT_3A55 16'h3946
`define CUBE_LUT_3A56 16'h3947
`define CUBE_LUT_3A57 16'h3947
`define CUBE_LUT_3A58 16'h3948
`define CUBE_LUT_3A59 16'h3948
`define CUBE_LUT_3A5A 16'h3949
`define CUBE_LUT_3A5B 16'h394A
`define CUBE_LUT_3A5C 16'h394A
`define CUBE_LUT_3A5D 16'h394B
`define CUBE_LUT_3A5E 16'h394B
`define CUBE_LUT_3A5F 16'h394C
`define CUBE_LUT_3A60 16'h394C
`define CUBE_LUT_3A61 16'h394D
`define CUBE_LUT_3A62 16'h394D
`define CUBE_LUT_3A63 16'h394E
`define CUBE_LUT_3A64 16'h394F
`define CUBE_LUT_3A65 16'h394F
`define CUBE_LUT_3A66 16'h3950
`define CUBE_LUT_3A67 16'h3950
`define CUBE_LUT_3A68 16'h3951
`define CUBE_LUT_3A69 16'h3951
`define CUBE_LUT_3A6A 16'h3952
`define CUBE_LUT_3A6B 16'h3953
`define CUBE_LUT_3A6C 16'h3953
`define CUBE_LUT_3A6D 16'h3954
`define CUBE_LUT_3A6E 16'h3954
`define CUBE_LUT_3A6F 16'h3955
`define CUBE_LUT_3A70 16'h3955
`define CUBE_LUT_3A71 16'h3956
`define CUBE_LUT_3A72 16'h3956
`define CUBE_LUT_3A73 16'h3957
`define CUBE_LUT_3A74 16'h3958
`define CUBE_LUT_3A75 16'h3958
`define CUBE_LUT_3A76 16'h3959
`define CUBE_LUT_3A77 16'h3959
`define CUBE_LUT_3A78 16'h395A
`define CUBE_LUT_3A79 16'h395A
`define CUBE_LUT_3A7A 16'h395B
`define CUBE_LUT_3A7B 16'h395B
`define CUBE_LUT_3A7C 16'h395C
`define CUBE_LUT_3A7D 16'h395C
`define CUBE_LUT_3A7E 16'h395D
`define CUBE_LUT_3A7F 16'h395E
`define CUBE_LUT_3A80 16'h395E
`define CUBE_LUT_3A81 16'h395F
`define CUBE_LUT_3A82 16'h395F
`define CUBE_LUT_3A83 16'h3960
`define CUBE_LUT_3A84 16'h3960
`define CUBE_LUT_3A85 16'h3961
`define CUBE_LUT_3A86 16'h3961
`define CUBE_LUT_3A87 16'h3962
`define CUBE_LUT_3A88 16'h3963
`define CUBE_LUT_3A89 16'h3963
`define CUBE_LUT_3A8A 16'h3964
`define CUBE_LUT_3A8B 16'h3964
`define CUBE_LUT_3A8C 16'h3965
`define CUBE_LUT_3A8D 16'h3965
`define CUBE_LUT_3A8E 16'h3966
`define CUBE_LUT_3A8F 16'h3966
`define CUBE_LUT_3A90 16'h3967
`define CUBE_LUT_3A91 16'h3967
`define CUBE_LUT_3A92 16'h3968
`define CUBE_LUT_3A93 16'h3969
`define CUBE_LUT_3A94 16'h3969
`define CUBE_LUT_3A95 16'h396A
`define CUBE_LUT_3A96 16'h396A
`define CUBE_LUT_3A97 16'h396B
`define CUBE_LUT_3A98 16'h396B
`define CUBE_LUT_3A99 16'h396C
`define CUBE_LUT_3A9A 16'h396C
`define CUBE_LUT_3A9B 16'h396D
`define CUBE_LUT_3A9C 16'h396D
`define CUBE_LUT_3A9D 16'h396E
`define CUBE_LUT_3A9E 16'h396E
`define CUBE_LUT_3A9F 16'h396F
`define CUBE_LUT_3AA0 16'h3970
`define CUBE_LUT_3AA1 16'h3970
`define CUBE_LUT_3AA2 16'h3971
`define CUBE_LUT_3AA3 16'h3971
`define CUBE_LUT_3AA4 16'h3972
`define CUBE_LUT_3AA5 16'h3972
`define CUBE_LUT_3AA6 16'h3973
`define CUBE_LUT_3AA7 16'h3973
`define CUBE_LUT_3AA8 16'h3974
`define CUBE_LUT_3AA9 16'h3974
`define CUBE_LUT_3AAA 16'h3975
`define CUBE_LUT_3AAB 16'h3975
`define CUBE_LUT_3AAC 16'h3976
`define CUBE_LUT_3AAD 16'h3977
`define CUBE_LUT_3AAE 16'h3977
`define CUBE_LUT_3AAF 16'h3978
`define CUBE_LUT_3AB0 16'h3978
`define CUBE_LUT_3AB1 16'h3979
`define CUBE_LUT_3AB2 16'h3979
`define CUBE_LUT_3AB3 16'h397A
`define CUBE_LUT_3AB4 16'h397A
`define CUBE_LUT_3AB5 16'h397B
`define CUBE_LUT_3AB6 16'h397B
`define CUBE_LUT_3AB7 16'h397C
`define CUBE_LUT_3AB8 16'h397C
`define CUBE_LUT_3AB9 16'h397D
`define CUBE_LUT_3ABA 16'h397D
`define CUBE_LUT_3ABB 16'h397E
`define CUBE_LUT_3ABC 16'h397E
`define CUBE_LUT_3ABD 16'h397F
`define CUBE_LUT_3ABE 16'h3980
`define CUBE_LUT_3ABF 16'h3980
`define CUBE_LUT_3AC0 16'h3981
`define CUBE_LUT_3AC1 16'h3981
`define CUBE_LUT_3AC2 16'h3982
`define CUBE_LUT_3AC3 16'h3982
`define CUBE_LUT_3AC4 16'h3983
`define CUBE_LUT_3AC5 16'h3983
`define CUBE_LUT_3AC6 16'h3984
`define CUBE_LUT_3AC7 16'h3984
`define CUBE_LUT_3AC8 16'h3985
`define CUBE_LUT_3AC9 16'h3985
`define CUBE_LUT_3ACA 16'h3986
`define CUBE_LUT_3ACB 16'h3986
`define CUBE_LUT_3ACC 16'h3987
`define CUBE_LUT_3ACD 16'h3987
`define CUBE_LUT_3ACE 16'h3988
`define CUBE_LUT_3ACF 16'h3988
`define CUBE_LUT_3AD0 16'h3989
`define CUBE_LUT_3AD1 16'h398A
`define CUBE_LUT_3AD2 16'h398A
`define CUBE_LUT_3AD3 16'h398B
`define CUBE_LUT_3AD4 16'h398B
`define CUBE_LUT_3AD5 16'h398C
`define CUBE_LUT_3AD6 16'h398C
`define CUBE_LUT_3AD7 16'h398D
`define CUBE_LUT_3AD8 16'h398D
`define CUBE_LUT_3AD9 16'h398E
`define CUBE_LUT_3ADA 16'h398E
`define CUBE_LUT_3ADB 16'h398F
`define CUBE_LUT_3ADC 16'h398F
`define CUBE_LUT_3ADD 16'h3990
`define CUBE_LUT_3ADE 16'h3990
`define CUBE_LUT_3ADF 16'h3991
`define CUBE_LUT_3AE0 16'h3991
`define CUBE_LUT_3AE1 16'h3992
`define CUBE_LUT_3AE2 16'h3992
`define CUBE_LUT_3AE3 16'h3993
`define CUBE_LUT_3AE4 16'h3993
`define CUBE_LUT_3AE5 16'h3994
`define CUBE_LUT_3AE6 16'h3994
`define CUBE_LUT_3AE7 16'h3995
`define CUBE_LUT_3AE8 16'h3995
`define CUBE_LUT_3AE9 16'h3996
`define CUBE_LUT_3AEA 16'h3996
`define CUBE_LUT_3AEB 16'h3997
`define CUBE_LUT_3AEC 16'h3997
`define CUBE_LUT_3AED 16'h3998
`define CUBE_LUT_3AEE 16'h3998
`define CUBE_LUT_3AEF 16'h3999
`define CUBE_LUT_3AF0 16'h3999
`define CUBE_LUT_3AF1 16'h399A
`define CUBE_LUT_3AF2 16'h399B
`define CUBE_LUT_3AF3 16'h399B
`define CUBE_LUT_3AF4 16'h399C
`define CUBE_LUT_3AF5 16'h399C
`define CUBE_LUT_3AF6 16'h399D
`define CUBE_LUT_3AF7 16'h399D
`define CUBE_LUT_3AF8 16'h399E
`define CUBE_LUT_3AF9 16'h399E
`define CUBE_LUT_3AFA 16'h399F
`define CUBE_LUT_3AFB 16'h399F
`define CUBE_LUT_3AFC 16'h39A0
`define CUBE_LUT_3AFD 16'h39A0
`define CUBE_LUT_3AFE 16'h39A1
`define CUBE_LUT_3AFF 16'h39A1
`define CUBE_LUT_3B00 16'h39A2
`define CUBE_LUT_3B01 16'h39A2
`define CUBE_LUT_3B02 16'h39A3
`define CUBE_LUT_3B03 16'h39A3
`define CUBE_LUT_3B04 16'h39A4
`define CUBE_LUT_3B05 16'h39A4
`define CUBE_LUT_3B06 16'h39A5
`define CUBE_LUT_3B07 16'h39A5
`define CUBE_LUT_3B08 16'h39A6
`define CUBE_LUT_3B09 16'h39A6
`define CUBE_LUT_3B0A 16'h39A7
`define CUBE_LUT_3B0B 16'h39A7
`define CUBE_LUT_3B0C 16'h39A8
`define CUBE_LUT_3B0D 16'h39A8
`define CUBE_LUT_3B0E 16'h39A9
`define CUBE_LUT_3B0F 16'h39A9
`define CUBE_LUT_3B10 16'h39AA
`define CUBE_LUT_3B11 16'h39AA
`define CUBE_LUT_3B12 16'h39AB
`define CUBE_LUT_3B13 16'h39AB
`define CUBE_LUT_3B14 16'h39AC
`define CUBE_LUT_3B15 16'h39AC
`define CUBE_LUT_3B16 16'h39AD
`define CUBE_LUT_3B17 16'h39AD
`define CUBE_LUT_3B18 16'h39AE
`define CUBE_LUT_3B19 16'h39AE
`define CUBE_LUT_3B1A 16'h39AF
`define CUBE_LUT_3B1B 16'h39AF
`define CUBE_LUT_3B1C 16'h39B0
`define CUBE_LUT_3B1D 16'h39B0
`define CUBE_LUT_3B1E 16'h39B1
`define CUBE_LUT_3B1F 16'h39B1
`define CUBE_LUT_3B20 16'h39B2
`define CUBE_LUT_3B21 16'h39B2
`define CUBE_LUT_3B22 16'h39B3
`define CUBE_LUT_3B23 16'h39B3
`define CUBE_LUT_3B24 16'h39B4
`define CUBE_LUT_3B25 16'h39B4
`define CUBE_LUT_3B26 16'h39B5
`define CUBE_LUT_3B27 16'h39B5
`define CUBE_LUT_3B28 16'h39B6
`define CUBE_LUT_3B29 16'h39B6
`define CUBE_LUT_3B2A 16'h39B6
`define CUBE_LUT_3B2B 16'h39B7
`define CUBE_LUT_3B2C 16'h39B7
`define CUBE_LUT_3B2D 16'h39B8
`define CUBE_LUT_3B2E 16'h39B8
`define CUBE_LUT_3B2F 16'h39B9
`define CUBE_LUT_3B30 16'h39B9
`define CUBE_LUT_3B31 16'h39BA
`define CUBE_LUT_3B32 16'h39BA
`define CUBE_LUT_3B33 16'h39BB
`define CUBE_LUT_3B34 16'h39BB
`define CUBE_LUT_3B35 16'h39BC
`define CUBE_LUT_3B36 16'h39BC
`define CUBE_LUT_3B37 16'h39BD
`define CUBE_LUT_3B38 16'h39BD
`define CUBE_LUT_3B39 16'h39BE
`define CUBE_LUT_3B3A 16'h39BE
`define CUBE_LUT_3B3B 16'h39BF
`define CUBE_LUT_3B3C 16'h39BF
`define CUBE_LUT_3B3D 16'h39C0
`define CUBE_LUT_3B3E 16'h39C0
`define CUBE_LUT_3B3F 16'h39C1
`define CUBE_LUT_3B40 16'h39C1
`define CUBE_LUT_3B41 16'h39C2
`define CUBE_LUT_3B42 16'h39C2
`define CUBE_LUT_3B43 16'h39C3
`define CUBE_LUT_3B44 16'h39C3
`define CUBE_LUT_3B45 16'h39C4
`define CUBE_LUT_3B46 16'h39C4
`define CUBE_LUT_3B47 16'h39C5
`define CUBE_LUT_3B48 16'h39C5
`define CUBE_LUT_3B49 16'h39C6
`define CUBE_LUT_3B4A 16'h39C6
`define CUBE_LUT_3B4B 16'h39C6
`define CUBE_LUT_3B4C 16'h39C7
`define CUBE_LUT_3B4D 16'h39C7
`define CUBE_LUT_3B4E 16'h39C8
`define CUBE_LUT_3B4F 16'h39C8
`define CUBE_LUT_3B50 16'h39C9
`define CUBE_LUT_3B51 16'h39C9
`define CUBE_LUT_3B52 16'h39CA
`define CUBE_LUT_3B53 16'h39CA
`define CUBE_LUT_3B54 16'h39CB
`define CUBE_LUT_3B55 16'h39CB
`define CUBE_LUT_3B56 16'h39CC
`define CUBE_LUT_3B57 16'h39CC
`define CUBE_LUT_3B58 16'h39CD
`define CUBE_LUT_3B59 16'h39CD
`define CUBE_LUT_3B5A 16'h39CE
`define CUBE_LUT_3B5B 16'h39CE
`define CUBE_LUT_3B5C 16'h39CF
`define CUBE_LUT_3B5D 16'h39CF
`define CUBE_LUT_3B5E 16'h39D0
`define CUBE_LUT_3B5F 16'h39D0
`define CUBE_LUT_3B60 16'h39D0
`define CUBE_LUT_3B61 16'h39D1
`define CUBE_LUT_3B62 16'h39D1
`define CUBE_LUT_3B63 16'h39D2
`define CUBE_LUT_3B64 16'h39D2
`define CUBE_LUT_3B65 16'h39D3
`define CUBE_LUT_3B66 16'h39D3
`define CUBE_LUT_3B67 16'h39D4
`define CUBE_LUT_3B68 16'h39D4
`define CUBE_LUT_3B69 16'h39D5
`define CUBE_LUT_3B6A 16'h39D5
`define CUBE_LUT_3B6B 16'h39D6
`define CUBE_LUT_3B6C 16'h39D6
`define CUBE_LUT_3B6D 16'h39D7
`define CUBE_LUT_3B6E 16'h39D7
`define CUBE_LUT_3B6F 16'h39D7
`define CUBE_LUT_3B70 16'h39D8
`define CUBE_LUT_3B71 16'h39D8
`define CUBE_LUT_3B72 16'h39D9
`define CUBE_LUT_3B73 16'h39D9
`define CUBE_LUT_3B74 16'h39DA
`define CUBE_LUT_3B75 16'h39DA
`define CUBE_LUT_3B76 16'h39DB
`define CUBE_LUT_3B77 16'h39DB
`define CUBE_LUT_3B78 16'h39DC
`define CUBE_LUT_3B79 16'h39DC
`define CUBE_LUT_3B7A 16'h39DD
`define CUBE_LUT_3B7B 16'h39DD
`define CUBE_LUT_3B7C 16'h39DE
`define CUBE_LUT_3B7D 16'h39DE
`define CUBE_LUT_3B7E 16'h39DE
`define CUBE_LUT_3B7F 16'h39DF
`define CUBE_LUT_3B80 16'h39DF
`define CUBE_LUT_3B81 16'h39E0
`define CUBE_LUT_3B82 16'h39E0
`define CUBE_LUT_3B83 16'h39E1
`define CUBE_LUT_3B84 16'h39E1
`define CUBE_LUT_3B85 16'h39E2
`define CUBE_LUT_3B86 16'h39E2
`define CUBE_LUT_3B87 16'h39E3
`define CUBE_LUT_3B88 16'h39E3
`define CUBE_LUT_3B89 16'h39E4
`define CUBE_LUT_3B8A 16'h39E4
`define CUBE_LUT_3B8B 16'h39E4
`define CUBE_LUT_3B8C 16'h39E5
`define CUBE_LUT_3B8D 16'h39E5
`define CUBE_LUT_3B8E 16'h39E6
`define CUBE_LUT_3B8F 16'h39E6
`define CUBE_LUT_3B90 16'h39E7
`define CUBE_LUT_3B91 16'h39E7
`define CUBE_LUT_3B92 16'h39E8
`define CUBE_LUT_3B93 16'h39E8
`define CUBE_LUT_3B94 16'h39E9
`define CUBE_LUT_3B95 16'h39E9
`define CUBE_LUT_3B96 16'h39E9
`define CUBE_LUT_3B97 16'h39EA
`define CUBE_LUT_3B98 16'h39EA
`define CUBE_LUT_3B99 16'h39EB
`define CUBE_LUT_3B9A 16'h39EB
`define CUBE_LUT_3B9B 16'h39EC
`define CUBE_LUT_3B9C 16'h39EC
`define CUBE_LUT_3B9D 16'h39ED
`define CUBE_LUT_3B9E 16'h39ED
`define CUBE_LUT_3B9F 16'h39EE
`define CUBE_LUT_3BA0 16'h39EE
`define CUBE_LUT_3BA1 16'h39EE
`define CUBE_LUT_3BA2 16'h39EF
`define CUBE_LUT_3BA3 16'h39EF
`define CUBE_LUT_3BA4 16'h39F0
`define CUBE_LUT_3BA5 16'h39F0
`define CUBE_LUT_3BA6 16'h39F1
`define CUBE_LUT_3BA7 16'h39F1
`define CUBE_LUT_3BA8 16'h39F2
`define CUBE_LUT_3BA9 16'h39F2
`define CUBE_LUT_3BAA 16'h39F2
`define CUBE_LUT_3BAB 16'h39F3
`define CUBE_LUT_3BAC 16'h39F3
`define CUBE_LUT_3BAD 16'h39F4
`define CUBE_LUT_3BAE 16'h39F4
`define CUBE_LUT_3BAF 16'h39F5
`define CUBE_LUT_3BB0 16'h39F5
`define CUBE_LUT_3BB1 16'h39F6
`define CUBE_LUT_3BB2 16'h39F6
`define CUBE_LUT_3BB3 16'h39F6
`define CUBE_LUT_3BB4 16'h39F7
`define CUBE_LUT_3BB5 16'h39F7
`define CUBE_LUT_3BB6 16'h39F8
`define CUBE_LUT_3BB7 16'h39F8
`define CUBE_LUT_3BB8 16'h39F9
`define CUBE_LUT_3BB9 16'h39F9
`define CUBE_LUT_3BBA 16'h39FA
`define CUBE_LUT_3BBB 16'h39FA
`define CUBE_LUT_3BBC 16'h39FA
`define CUBE_LUT_3BBD 16'h39FB
`define CUBE_LUT_3BBE 16'h39FB
`define CUBE_LUT_3BBF 16'h39FC
`define CUBE_LUT_3BC0 16'h39FC
`define CUBE_LUT_3BC1 16'h39FD
`define CUBE_LUT_3BC2 16'h39FD
`define CUBE_LUT_3BC3 16'h39FE
`define CUBE_LUT_3BC4 16'h39FE
`define CUBE_LUT_3BC5 16'h39FE
`define CUBE_LUT_3BC6 16'h39FF
`define CUBE_LUT_3BC7 16'h39FF
`define CUBE_LUT_3BC8 16'h3A00
`define CUBE_LUT_3BC9 16'h3A00
`define CUBE_LUT_3BCA 16'h3A01
`define CUBE_LUT_3BCB 16'h3A01
`define CUBE_LUT_3BCC 16'h3A01
`define CUBE_LUT_3BCD 16'h3A02
`define CUBE_LUT_3BCE 16'h3A02
`define CUBE_LUT_3BCF 16'h3A03
`define CUBE_LUT_3BD0 16'h3A03
`define CUBE_LUT_3BD1 16'h3A04
`define CUBE_LUT_3BD2 16'h3A04
`define CUBE_LUT_3BD3 16'h3A05
`define CUBE_LUT_3BD4 16'h3A05
`define CUBE_LUT_3BD5 16'h3A05
`define CUBE_LUT_3BD6 16'h3A06
`define CUBE_LUT_3BD7 16'h3A06
`define CUBE_LUT_3BD8 16'h3A07
`define CUBE_LUT_3BD9 16'h3A07
`define CUBE_LUT_3BDA 16'h3A08
`define CUBE_LUT_3BDB 16'h3A08
`define CUBE_LUT_3BDC 16'h3A08
`define CUBE_LUT_3BDD 16'h3A09
`define CUBE_LUT_3BDE 16'h3A09
`define CUBE_LUT_3BDF 16'h3A0A
`define CUBE_LUT_3BE0 16'h3A0A
`define CUBE_LUT_3BE1 16'h3A0B
`define CUBE_LUT_3BE2 16'h3A0B
`define CUBE_LUT_3BE3 16'h3A0B
`define CUBE_LUT_3BE4 16'h3A0C
`define CUBE_LUT_3BE5 16'h3A0C
`define CUBE_LUT_3BE6 16'h3A0D
`define CUBE_LUT_3BE7 16'h3A0D
`define CUBE_LUT_3BE8 16'h3A0E
`define CUBE_LUT_3BE9 16'h3A0E
`define CUBE_LUT_3BEA 16'h3A0E
`define CUBE_LUT_3BEB 16'h3A0F
`define CUBE_LUT_3BEC 16'h3A0F
`define CUBE_LUT_3BED 16'h3A10
`define CUBE_LUT_3BEE 16'h3A10
`define CUBE_LUT_3BEF 16'h3A11
`define CUBE_LUT_3BF0 16'h3A11
`define CUBE_LUT_3BF1 16'h3A11
`define CUBE_LUT_3BF2 16'h3A12
`define CUBE_LUT_3BF3 16'h3A12
`define CUBE_LUT_3BF4 16'h3A13
`define CUBE_LUT_3BF5 16'h3A13
`define CUBE_LUT_3BF6 16'h3A14
`define CUBE_LUT_3BF7 16'h3A14
`define CUBE_LUT_3BF8 16'h3A14
`define CUBE_LUT_3BF9 16'h3A15
`define CUBE_LUT_3BFA 16'h3A15
`define CUBE_LUT_3BFB 16'h3A16
`define CUBE_LUT_3BFC 16'h3A16
`define CUBE_LUT_3BFD 16'h3A16
`define CUBE_LUT_3BFE 16'h3A17
`define CUBE_LUT_3BFF 16'h3A17
`define CUBE_LUT_3C00 16'h3A18
`define CUBE_LUT_3C01 16'h3A19
`define CUBE_LUT_3C02 16'h3A19
`define CUBE_LUT_3C03 16'h3A1A
`define CUBE_LUT_3C04 16'h3A1B
`define CUBE_LUT_3C05 16'h3A1C
`define CUBE_LUT_3C06 16'h3A1D
`define CUBE_LUT_3C07 16'h3A1E
`define CUBE_LUT_3C08 16'h3A1E
`define CUBE_LUT_3C09 16'h3A1F
`define CUBE_LUT_3C0A 16'h3A20
`define CUBE_LUT_3C0B 16'h3A21
`define CUBE_LUT_3C0C 16'h3A22
`define CUBE_LUT_3C0D 16'h3A23
`define CUBE_LUT_3C0E 16'h3A23
`define CUBE_LUT_3C0F 16'h3A24
`define CUBE_LUT_3C10 16'h3A25
`define CUBE_LUT_3C11 16'h3A26
`define CUBE_LUT_3C12 16'h3A27
`define CUBE_LUT_3C13 16'h3A27
`define CUBE_LUT_3C14 16'h3A28
`define CUBE_LUT_3C15 16'h3A29
`define CUBE_LUT_3C16 16'h3A2A
`define CUBE_LUT_3C17 16'h3A2B
`define CUBE_LUT_3C18 16'h3A2C
`define CUBE_LUT_3C19 16'h3A2C
`define CUBE_LUT_3C1A 16'h3A2D
`define CUBE_LUT_3C1B 16'h3A2E
`define CUBE_LUT_3C1C 16'h3A2F
`define CUBE_LUT_3C1D 16'h3A30
`define CUBE_LUT_3C1E 16'h3A30
`define CUBE_LUT_3C1F 16'h3A31
`define CUBE_LUT_3C20 16'h3A32
`define CUBE_LUT_3C21 16'h3A33
`define CUBE_LUT_3C22 16'h3A34
`define CUBE_LUT_3C23 16'h3A34
`define CUBE_LUT_3C24 16'h3A35
`define CUBE_LUT_3C25 16'h3A36
`define CUBE_LUT_3C26 16'h3A37
`define CUBE_LUT_3C27 16'h3A38
`define CUBE_LUT_3C28 16'h3A38
`define CUBE_LUT_3C29 16'h3A39
`define CUBE_LUT_3C2A 16'h3A3A
`define CUBE_LUT_3C2B 16'h3A3B
`define CUBE_LUT_3C2C 16'h3A3C
`define CUBE_LUT_3C2D 16'h3A3C
`define CUBE_LUT_3C2E 16'h3A3D
`define CUBE_LUT_3C2F 16'h3A3E
`define CUBE_LUT_3C30 16'h3A3F
`define CUBE_LUT_3C31 16'h3A3F
`define CUBE_LUT_3C32 16'h3A40
`define CUBE_LUT_3C33 16'h3A41
`define CUBE_LUT_3C34 16'h3A42
`define CUBE_LUT_3C35 16'h3A43
`define CUBE_LUT_3C36 16'h3A43
`define CUBE_LUT_3C37 16'h3A44
`define CUBE_LUT_3C38 16'h3A45
`define CUBE_LUT_3C39 16'h3A46
`define CUBE_LUT_3C3A 16'h3A46
`define CUBE_LUT_3C3B 16'h3A47
`define CUBE_LUT_3C3C 16'h3A48
`define CUBE_LUT_3C3D 16'h3A49
`define CUBE_LUT_3C3E 16'h3A49
`define CUBE_LUT_3C3F 16'h3A4A
`define CUBE_LUT_3C40 16'h3A4B
`define CUBE_LUT_3C41 16'h3A4C
`define CUBE_LUT_3C42 16'h3A4D
`define CUBE_LUT_3C43 16'h3A4D
`define CUBE_LUT_3C44 16'h3A4E
`define CUBE_LUT_3C45 16'h3A4F
`define CUBE_LUT_3C46 16'h3A50
`define CUBE_LUT_3C47 16'h3A50
`define CUBE_LUT_3C48 16'h3A51
`define CUBE_LUT_3C49 16'h3A52
`define CUBE_LUT_3C4A 16'h3A53
`define CUBE_LUT_3C4B 16'h3A53
`define CUBE_LUT_3C4C 16'h3A54
`define CUBE_LUT_3C4D 16'h3A55
`define CUBE_LUT_3C4E 16'h3A56
`define CUBE_LUT_3C4F 16'h3A56
`define CUBE_LUT_3C50 16'h3A57
`define CUBE_LUT_3C51 16'h3A58
`define CUBE_LUT_3C52 16'h3A59
`define CUBE_LUT_3C53 16'h3A59
`define CUBE_LUT_3C54 16'h3A5A
`define CUBE_LUT_3C55 16'h3A5B
`define CUBE_LUT_3C56 16'h3A5B
`define CUBE_LUT_3C57 16'h3A5C
`define CUBE_LUT_3C58 16'h3A5D
`define CUBE_LUT_3C59 16'h3A5E
`define CUBE_LUT_3C5A 16'h3A5E
`define CUBE_LUT_3C5B 16'h3A5F
`define CUBE_LUT_3C5C 16'h3A60
`define CUBE_LUT_3C5D 16'h3A61
`define CUBE_LUT_3C5E 16'h3A61
`define CUBE_LUT_3C5F 16'h3A62
`define CUBE_LUT_3C60 16'h3A63
`define CUBE_LUT_3C61 16'h3A64
`define CUBE_LUT_3C62 16'h3A64
`define CUBE_LUT_3C63 16'h3A65
`define CUBE_LUT_3C64 16'h3A66
`define CUBE_LUT_3C65 16'h3A66
`define CUBE_LUT_3C66 16'h3A67
`define CUBE_LUT_3C67 16'h3A68
`define CUBE_LUT_3C68 16'h3A69
`define CUBE_LUT_3C69 16'h3A69
`define CUBE_LUT_3C6A 16'h3A6A
`define CUBE_LUT_3C6B 16'h3A6B
`define CUBE_LUT_3C6C 16'h3A6B
`define CUBE_LUT_3C6D 16'h3A6C
`define CUBE_LUT_3C6E 16'h3A6D
`define CUBE_LUT_3C6F 16'h3A6E
`define CUBE_LUT_3C70 16'h3A6E
`define CUBE_LUT_3C71 16'h3A6F
`define CUBE_LUT_3C72 16'h3A70
`define CUBE_LUT_3C73 16'h3A70
`define CUBE_LUT_3C74 16'h3A71
`define CUBE_LUT_3C75 16'h3A72
`define CUBE_LUT_3C76 16'h3A72
`define CUBE_LUT_3C77 16'h3A73
`define CUBE_LUT_3C78 16'h3A74
`define CUBE_LUT_3C79 16'h3A75
`define CUBE_LUT_3C7A 16'h3A75
`define CUBE_LUT_3C7B 16'h3A76
`define CUBE_LUT_3C7C 16'h3A77
`define CUBE_LUT_3C7D 16'h3A77
`define CUBE_LUT_3C7E 16'h3A78
`define CUBE_LUT_3C7F 16'h3A79
`define CUBE_LUT_3C80 16'h3A79
`define CUBE_LUT_3C81 16'h3A7A
`define CUBE_LUT_3C82 16'h3A7B
`define CUBE_LUT_3C83 16'h3A7C
`define CUBE_LUT_3C84 16'h3A7C
`define CUBE_LUT_3C85 16'h3A7D
`define CUBE_LUT_3C86 16'h3A7E
`define CUBE_LUT_3C87 16'h3A7E
`define CUBE_LUT_3C88 16'h3A7F
`define CUBE_LUT_3C89 16'h3A80
`define CUBE_LUT_3C8A 16'h3A80
`define CUBE_LUT_3C8B 16'h3A81
`define CUBE_LUT_3C8C 16'h3A82
`define CUBE_LUT_3C8D 16'h3A82
`define CUBE_LUT_3C8E 16'h3A83
`define CUBE_LUT_3C8F 16'h3A84
`define CUBE_LUT_3C90 16'h3A84
`define CUBE_LUT_3C91 16'h3A85
`define CUBE_LUT_3C92 16'h3A86
`define CUBE_LUT_3C93 16'h3A86
`define CUBE_LUT_3C94 16'h3A87
`define CUBE_LUT_3C95 16'h3A88
`define CUBE_LUT_3C96 16'h3A88
`define CUBE_LUT_3C97 16'h3A89
`define CUBE_LUT_3C98 16'h3A8A
`define CUBE_LUT_3C99 16'h3A8A
`define CUBE_LUT_3C9A 16'h3A8B
`define CUBE_LUT_3C9B 16'h3A8C
`define CUBE_LUT_3C9C 16'h3A8C
`define CUBE_LUT_3C9D 16'h3A8D
`define CUBE_LUT_3C9E 16'h3A8E
`define CUBE_LUT_3C9F 16'h3A8E
`define CUBE_LUT_3CA0 16'h3A8F
`define CUBE_LUT_3CA1 16'h3A90
`define CUBE_LUT_3CA2 16'h3A90
`define CUBE_LUT_3CA3 16'h3A91
`define CUBE_LUT_3CA4 16'h3A92
`define CUBE_LUT_3CA5 16'h3A92
`define CUBE_LUT_3CA6 16'h3A93
`define CUBE_LUT_3CA7 16'h3A94
`define CUBE_LUT_3CA8 16'h3A94
`define CUBE_LUT_3CA9 16'h3A95
`define CUBE_LUT_3CAA 16'h3A95
`define CUBE_LUT_3CAB 16'h3A96
`define CUBE_LUT_3CAC 16'h3A97
`define CUBE_LUT_3CAD 16'h3A97
`define CUBE_LUT_3CAE 16'h3A98
`define CUBE_LUT_3CAF 16'h3A99
`define CUBE_LUT_3CB0 16'h3A99
`define CUBE_LUT_3CB1 16'h3A9A
`define CUBE_LUT_3CB2 16'h3A9B
`define CUBE_LUT_3CB3 16'h3A9B
`define CUBE_LUT_3CB4 16'h3A9C
`define CUBE_LUT_3CB5 16'h3A9D
`define CUBE_LUT_3CB6 16'h3A9D
`define CUBE_LUT_3CB7 16'h3A9E
`define CUBE_LUT_3CB8 16'h3A9E
`define CUBE_LUT_3CB9 16'h3A9F
`define CUBE_LUT_3CBA 16'h3AA0
`define CUBE_LUT_3CBB 16'h3AA0
`define CUBE_LUT_3CBC 16'h3AA1
`define CUBE_LUT_3CBD 16'h3AA2
`define CUBE_LUT_3CBE 16'h3AA2
`define CUBE_LUT_3CBF 16'h3AA3
`define CUBE_LUT_3CC0 16'h3AA3
`define CUBE_LUT_3CC1 16'h3AA4
`define CUBE_LUT_3CC2 16'h3AA5
`define CUBE_LUT_3CC3 16'h3AA5
`define CUBE_LUT_3CC4 16'h3AA6
`define CUBE_LUT_3CC5 16'h3AA7
`define CUBE_LUT_3CC6 16'h3AA7
`define CUBE_LUT_3CC7 16'h3AA8
`define CUBE_LUT_3CC8 16'h3AA8
`define CUBE_LUT_3CC9 16'h3AA9
`define CUBE_LUT_3CCA 16'h3AAA
`define CUBE_LUT_3CCB 16'h3AAA
`define CUBE_LUT_3CCC 16'h3AAB
`define CUBE_LUT_3CCD 16'h3AAB
`define CUBE_LUT_3CCE 16'h3AAC
`define CUBE_LUT_3CCF 16'h3AAD
`define CUBE_LUT_3CD0 16'h3AAD
`define CUBE_LUT_3CD1 16'h3AAE
`define CUBE_LUT_3CD2 16'h3AAE
`define CUBE_LUT_3CD3 16'h3AAF
`define CUBE_LUT_3CD4 16'h3AB0
`define CUBE_LUT_3CD5 16'h3AB0
`define CUBE_LUT_3CD6 16'h3AB1
`define CUBE_LUT_3CD7 16'h3AB1
`define CUBE_LUT_3CD8 16'h3AB2
`define CUBE_LUT_3CD9 16'h3AB3
`define CUBE_LUT_3CDA 16'h3AB3
`define CUBE_LUT_3CDB 16'h3AB4
`define CUBE_LUT_3CDC 16'h3AB4
`define CUBE_LUT_3CDD 16'h3AB5
`define CUBE_LUT_3CDE 16'h3AB6
`define CUBE_LUT_3CDF 16'h3AB6
`define CUBE_LUT_3CE0 16'h3AB7
`define CUBE_LUT_3CE1 16'h3AB7
`define CUBE_LUT_3CE2 16'h3AB8
`define CUBE_LUT_3CE3 16'h3AB9
`define CUBE_LUT_3CE4 16'h3AB9
`define CUBE_LUT_3CE5 16'h3ABA
`define CUBE_LUT_3CE6 16'h3ABA
`define CUBE_LUT_3CE7 16'h3ABB
`define CUBE_LUT_3CE8 16'h3ABC
`define CUBE_LUT_3CE9 16'h3ABC
`define CUBE_LUT_3CEA 16'h3ABD
`define CUBE_LUT_3CEB 16'h3ABD
`define CUBE_LUT_3CEC 16'h3ABE
`define CUBE_LUT_3CED 16'h3ABE
`define CUBE_LUT_3CEE 16'h3ABF
`define CUBE_LUT_3CEF 16'h3AC0
`define CUBE_LUT_3CF0 16'h3AC0
`define CUBE_LUT_3CF1 16'h3AC1
`define CUBE_LUT_3CF2 16'h3AC1
`define CUBE_LUT_3CF3 16'h3AC2
`define CUBE_LUT_3CF4 16'h3AC2
`define CUBE_LUT_3CF5 16'h3AC3
`define CUBE_LUT_3CF6 16'h3AC4
`define CUBE_LUT_3CF7 16'h3AC4
`define CUBE_LUT_3CF8 16'h3AC5
`define CUBE_LUT_3CF9 16'h3AC5
`define CUBE_LUT_3CFA 16'h3AC6
`define CUBE_LUT_3CFB 16'h3AC6
`define CUBE_LUT_3CFC 16'h3AC7
`define CUBE_LUT_3CFD 16'h3AC8
`define CUBE_LUT_3CFE 16'h3AC8
`define CUBE_LUT_3CFF 16'h3AC9
`define CUBE_LUT_3D00 16'h3AC9
`define CUBE_LUT_3D01 16'h3ACA
`define CUBE_LUT_3D02 16'h3ACA
`define CUBE_LUT_3D03 16'h3ACB
`define CUBE_LUT_3D04 16'h3ACC
`define CUBE_LUT_3D05 16'h3ACC
`define CUBE_LUT_3D06 16'h3ACD
`define CUBE_LUT_3D07 16'h3ACD
`define CUBE_LUT_3D08 16'h3ACE
`define CUBE_LUT_3D09 16'h3ACE
`define CUBE_LUT_3D0A 16'h3ACF
`define CUBE_LUT_3D0B 16'h3ACF
`define CUBE_LUT_3D0C 16'h3AD0
`define CUBE_LUT_3D0D 16'h3AD0
`define CUBE_LUT_3D0E 16'h3AD1
`define CUBE_LUT_3D0F 16'h3AD2
`define CUBE_LUT_3D10 16'h3AD2
`define CUBE_LUT_3D11 16'h3AD3
`define CUBE_LUT_3D12 16'h3AD3
`define CUBE_LUT_3D13 16'h3AD4
`define CUBE_LUT_3D14 16'h3AD4
`define CUBE_LUT_3D15 16'h3AD5
`define CUBE_LUT_3D16 16'h3AD5
`define CUBE_LUT_3D17 16'h3AD6
`define CUBE_LUT_3D18 16'h3AD6
`define CUBE_LUT_3D19 16'h3AD7
`define CUBE_LUT_3D1A 16'h3AD8
`define CUBE_LUT_3D1B 16'h3AD8
`define CUBE_LUT_3D1C 16'h3AD9
`define CUBE_LUT_3D1D 16'h3AD9
`define CUBE_LUT_3D1E 16'h3ADA
`define CUBE_LUT_3D1F 16'h3ADA
`define CUBE_LUT_3D20 16'h3ADB
`define CUBE_LUT_3D21 16'h3ADB
`define CUBE_LUT_3D22 16'h3ADC
`define CUBE_LUT_3D23 16'h3ADC
`define CUBE_LUT_3D24 16'h3ADD
`define CUBE_LUT_3D25 16'h3ADD
`define CUBE_LUT_3D26 16'h3ADE
`define CUBE_LUT_3D27 16'h3ADE
`define CUBE_LUT_3D28 16'h3ADF
`define CUBE_LUT_3D29 16'h3AE0
`define CUBE_LUT_3D2A 16'h3AE0
`define CUBE_LUT_3D2B 16'h3AE1
`define CUBE_LUT_3D2C 16'h3AE1
`define CUBE_LUT_3D2D 16'h3AE2
`define CUBE_LUT_3D2E 16'h3AE2
`define CUBE_LUT_3D2F 16'h3AE3
`define CUBE_LUT_3D30 16'h3AE3
`define CUBE_LUT_3D31 16'h3AE4
`define CUBE_LUT_3D32 16'h3AE4
`define CUBE_LUT_3D33 16'h3AE5
`define CUBE_LUT_3D34 16'h3AE5
`define CUBE_LUT_3D35 16'h3AE6
`define CUBE_LUT_3D36 16'h3AE6
`define CUBE_LUT_3D37 16'h3AE7
`define CUBE_LUT_3D38 16'h3AE7
`define CUBE_LUT_3D39 16'h3AE8
`define CUBE_LUT_3D3A 16'h3AE8
`define CUBE_LUT_3D3B 16'h3AE9
`define CUBE_LUT_3D3C 16'h3AE9
`define CUBE_LUT_3D3D 16'h3AEA
`define CUBE_LUT_3D3E 16'h3AEA
`define CUBE_LUT_3D3F 16'h3AEB
`define CUBE_LUT_3D40 16'h3AEB
`define CUBE_LUT_3D41 16'h3AEC
`define CUBE_LUT_3D42 16'h3AEC
`define CUBE_LUT_3D43 16'h3AED
`define CUBE_LUT_3D44 16'h3AED
`define CUBE_LUT_3D45 16'h3AEE
`define CUBE_LUT_3D46 16'h3AEE
`define CUBE_LUT_3D47 16'h3AEF
`define CUBE_LUT_3D48 16'h3AEF
`define CUBE_LUT_3D49 16'h3AF0
`define CUBE_LUT_3D4A 16'h3AF0
`define CUBE_LUT_3D4B 16'h3AF1
`define CUBE_LUT_3D4C 16'h3AF1
`define CUBE_LUT_3D4D 16'h3AF2
`define CUBE_LUT_3D4E 16'h3AF2
`define CUBE_LUT_3D4F 16'h3AF3
`define CUBE_LUT_3D50 16'h3AF3
`define CUBE_LUT_3D51 16'h3AF4
`define CUBE_LUT_3D52 16'h3AF4
`define CUBE_LUT_3D53 16'h3AF5
`define CUBE_LUT_3D54 16'h3AF5
`define CUBE_LUT_3D55 16'h3AF6
`define CUBE_LUT_3D56 16'h3AF6
`define CUBE_LUT_3D57 16'h3AF7
`define CUBE_LUT_3D58 16'h3AF7
`define CUBE_LUT_3D59 16'h3AF8
`define CUBE_LUT_3D5A 16'h3AF8
`define CUBE_LUT_3D5B 16'h3AF9
`define CUBE_LUT_3D5C 16'h3AF9
`define CUBE_LUT_3D5D 16'h3AFA
`define CUBE_LUT_3D5E 16'h3AFA
`define CUBE_LUT_3D5F 16'h3AFB
`define CUBE_LUT_3D60 16'h3AFB
`define CUBE_LUT_3D61 16'h3AFC
`define CUBE_LUT_3D62 16'h3AFC
`define CUBE_LUT_3D63 16'h3AFC
`define CUBE_LUT_3D64 16'h3AFD
`define CUBE_LUT_3D65 16'h3AFD
`define CUBE_LUT_3D66 16'h3AFE
`define CUBE_LUT_3D67 16'h3AFE
`define CUBE_LUT_3D68 16'h3AFF
`define CUBE_LUT_3D69 16'h3AFF
`define CUBE_LUT_3D6A 16'h3B00
`define CUBE_LUT_3D6B 16'h3B00
`define CUBE_LUT_3D6C 16'h3B01
`define CUBE_LUT_3D6D 16'h3B01
`define CUBE_LUT_3D6E 16'h3B02
`define CUBE_LUT_3D6F 16'h3B02
`define CUBE_LUT_3D70 16'h3B03
`define CUBE_LUT_3D71 16'h3B03
`define CUBE_LUT_3D72 16'h3B03
`define CUBE_LUT_3D73 16'h3B04
`define CUBE_LUT_3D74 16'h3B04
`define CUBE_LUT_3D75 16'h3B05
`define CUBE_LUT_3D76 16'h3B05
`define CUBE_LUT_3D77 16'h3B06
`define CUBE_LUT_3D78 16'h3B06
`define CUBE_LUT_3D79 16'h3B07
`define CUBE_LUT_3D7A 16'h3B07
`define CUBE_LUT_3D7B 16'h3B08
`define CUBE_LUT_3D7C 16'h3B08
`define CUBE_LUT_3D7D 16'h3B09
`define CUBE_LUT_3D7E 16'h3B09
`define CUBE_LUT_3D7F 16'h3B09
`define CUBE_LUT_3D80 16'h3B0A
`define CUBE_LUT_3D81 16'h3B0A
`define CUBE_LUT_3D82 16'h3B0B
`define CUBE_LUT_3D83 16'h3B0B
`define CUBE_LUT_3D84 16'h3B0C
`define CUBE_LUT_3D85 16'h3B0C
`define CUBE_LUT_3D86 16'h3B0D
`define CUBE_LUT_3D87 16'h3B0D
`define CUBE_LUT_3D88 16'h3B0D
`define CUBE_LUT_3D89 16'h3B0E
`define CUBE_LUT_3D8A 16'h3B0E
`define CUBE_LUT_3D8B 16'h3B0F
`define CUBE_LUT_3D8C 16'h3B0F
`define CUBE_LUT_3D8D 16'h3B10
`define CUBE_LUT_3D8E 16'h3B10
`define CUBE_LUT_3D8F 16'h3B11
`define CUBE_LUT_3D90 16'h3B11
`define CUBE_LUT_3D91 16'h3B11
`define CUBE_LUT_3D92 16'h3B12
`define CUBE_LUT_3D93 16'h3B12
`define CUBE_LUT_3D94 16'h3B13
`define CUBE_LUT_3D95 16'h3B13
`define CUBE_LUT_3D96 16'h3B14
`define CUBE_LUT_3D97 16'h3B14
`define CUBE_LUT_3D98 16'h3B15
`define CUBE_LUT_3D99 16'h3B15
`define CUBE_LUT_3D9A 16'h3B15
`define CUBE_LUT_3D9B 16'h3B16
`define CUBE_LUT_3D9C 16'h3B16
`define CUBE_LUT_3D9D 16'h3B17
`define CUBE_LUT_3D9E 16'h3B17
`define CUBE_LUT_3D9F 16'h3B18
`define CUBE_LUT_3DA0 16'h3B18
`define CUBE_LUT_3DA1 16'h3B18
`define CUBE_LUT_3DA2 16'h3B19
`define CUBE_LUT_3DA3 16'h3B19
`define CUBE_LUT_3DA4 16'h3B1A
`define CUBE_LUT_3DA5 16'h3B1A
`define CUBE_LUT_3DA6 16'h3B1B
`define CUBE_LUT_3DA7 16'h3B1B
`define CUBE_LUT_3DA8 16'h3B1B
`define CUBE_LUT_3DA9 16'h3B1C
`define CUBE_LUT_3DAA 16'h3B1C
`define CUBE_LUT_3DAB 16'h3B1D
`define CUBE_LUT_3DAC 16'h3B1D
`define CUBE_LUT_3DAD 16'h3B1D
`define CUBE_LUT_3DAE 16'h3B1E
`define CUBE_LUT_3DAF 16'h3B1E
`define CUBE_LUT_3DB0 16'h3B1F
`define CUBE_LUT_3DB1 16'h3B1F
`define CUBE_LUT_3DB2 16'h3B20
`define CUBE_LUT_3DB3 16'h3B20
`define CUBE_LUT_3DB4 16'h3B20
`define CUBE_LUT_3DB5 16'h3B21
`define CUBE_LUT_3DB6 16'h3B21
`define CUBE_LUT_3DB7 16'h3B22
`define CUBE_LUT_3DB8 16'h3B22
`define CUBE_LUT_3DB9 16'h3B22
`define CUBE_LUT_3DBA 16'h3B23
`define CUBE_LUT_3DBB 16'h3B23
`define CUBE_LUT_3DBC 16'h3B24
`define CUBE_LUT_3DBD 16'h3B24
`define CUBE_LUT_3DBE 16'h3B24
`define CUBE_LUT_3DBF 16'h3B25
`define CUBE_LUT_3DC0 16'h3B25
`define CUBE_LUT_3DC1 16'h3B26
`define CUBE_LUT_3DC2 16'h3B26
`define CUBE_LUT_3DC3 16'h3B26
`define CUBE_LUT_3DC4 16'h3B27
`define CUBE_LUT_3DC5 16'h3B27
`define CUBE_LUT_3DC6 16'h3B28
`define CUBE_LUT_3DC7 16'h3B28
`define CUBE_LUT_3DC8 16'h3B28
`define CUBE_LUT_3DC9 16'h3B29
`define CUBE_LUT_3DCA 16'h3B29
`define CUBE_LUT_3DCB 16'h3B2A
`define CUBE_LUT_3DCC 16'h3B2A
`define CUBE_LUT_3DCD 16'h3B2A
`define CUBE_LUT_3DCE 16'h3B2B
`define CUBE_LUT_3DCF 16'h3B2B
`define CUBE_LUT_3DD0 16'h3B2C
`define CUBE_LUT_3DD1 16'h3B2C
`define CUBE_LUT_3DD2 16'h3B2C
`define CUBE_LUT_3DD3 16'h3B2D
`define CUBE_LUT_3DD4 16'h3B2D
`define CUBE_LUT_3DD5 16'h3B2E
`define CUBE_LUT_3DD6 16'h3B2E
`define CUBE_LUT_3DD7 16'h3B2E
`define CUBE_LUT_3DD8 16'h3B2F
`define CUBE_LUT_3DD9 16'h3B2F
`define CUBE_LUT_3DDA 16'h3B30
`define CUBE_LUT_3DDB 16'h3B30
`define CUBE_LUT_3DDC 16'h3B30
`define CUBE_LUT_3DDD 16'h3B31
`define CUBE_LUT_3DDE 16'h3B31
`define CUBE_LUT_3DDF 16'h3B31
`define CUBE_LUT_3DE0 16'h3B32
`define CUBE_LUT_3DE1 16'h3B32
`define CUBE_LUT_3DE2 16'h3B33
`define CUBE_LUT_3DE3 16'h3B33
`define CUBE_LUT_3DE4 16'h3B33
`define CUBE_LUT_3DE5 16'h3B34
`define CUBE_LUT_3DE6 16'h3B34
`define CUBE_LUT_3DE7 16'h3B35
`define CUBE_LUT_3DE8 16'h3B35
`define CUBE_LUT_3DE9 16'h3B35
`define CUBE_LUT_3DEA 16'h3B36
`define CUBE_LUT_3DEB 16'h3B36
`define CUBE_LUT_3DEC 16'h3B36
`define CUBE_LUT_3DED 16'h3B37
`define CUBE_LUT_3DEE 16'h3B37
`define CUBE_LUT_3DEF 16'h3B38
`define CUBE_LUT_3DF0 16'h3B38
`define CUBE_LUT_3DF1 16'h3B38
`define CUBE_LUT_3DF2 16'h3B39
`define CUBE_LUT_3DF3 16'h3B39
`define CUBE_LUT_3DF4 16'h3B39
`define CUBE_LUT_3DF5 16'h3B3A
`define CUBE_LUT_3DF6 16'h3B3A
`define CUBE_LUT_3DF7 16'h3B3A
`define CUBE_LUT_3DF8 16'h3B3B
`define CUBE_LUT_3DF9 16'h3B3B
`define CUBE_LUT_3DFA 16'h3B3C
`define CUBE_LUT_3DFB 16'h3B3C
`define CUBE_LUT_3DFC 16'h3B3C
`define CUBE_LUT_3DFD 16'h3B3D
`define CUBE_LUT_3DFE 16'h3B3D
`define CUBE_LUT_3DFF 16'h3B3D
`define CUBE_LUT_3E00 16'h3B3E
`define CUBE_LUT_3E01 16'h3B3E
`define CUBE_LUT_3E02 16'h3B3E
`define CUBE_LUT_3E03 16'h3B3F
`define CUBE_LUT_3E04 16'h3B3F
`define CUBE_LUT_3E05 16'h3B40
`define CUBE_LUT_3E06 16'h3B40
`define CUBE_LUT_3E07 16'h3B40
`define CUBE_LUT_3E08 16'h3B41
`define CUBE_LUT_3E09 16'h3B41
`define CUBE_LUT_3E0A 16'h3B41
`define CUBE_LUT_3E0B 16'h3B42
`define CUBE_LUT_3E0C 16'h3B42
`define CUBE_LUT_3E0D 16'h3B42
`define CUBE_LUT_3E0E 16'h3B43
`define CUBE_LUT_3E0F 16'h3B43
`define CUBE_LUT_3E10 16'h3B43
`define CUBE_LUT_3E11 16'h3B44
`define CUBE_LUT_3E12 16'h3B44
`define CUBE_LUT_3E13 16'h3B44
`define CUBE_LUT_3E14 16'h3B45
`define CUBE_LUT_3E15 16'h3B45
`define CUBE_LUT_3E16 16'h3B46
`define CUBE_LUT_3E17 16'h3B46
`define CUBE_LUT_3E18 16'h3B46
`define CUBE_LUT_3E19 16'h3B47
`define CUBE_LUT_3E1A 16'h3B47
`define CUBE_LUT_3E1B 16'h3B47
`define CUBE_LUT_3E1C 16'h3B48
`define CUBE_LUT_3E1D 16'h3B48
`define CUBE_LUT_3E1E 16'h3B48
`define CUBE_LUT_3E1F 16'h3B49
`define CUBE_LUT_3E20 16'h3B49
`define CUBE_LUT_3E21 16'h3B49
`define CUBE_LUT_3E22 16'h3B4A
`define CUBE_LUT_3E23 16'h3B4A
`define CUBE_LUT_3E24 16'h3B4A
`define CUBE_LUT_3E25 16'h3B4B
`define CUBE_LUT_3E26 16'h3B4B
`define CUBE_LUT_3E27 16'h3B4B
`define CUBE_LUT_3E28 16'h3B4C
`define CUBE_LUT_3E29 16'h3B4C
`define CUBE_LUT_3E2A 16'h3B4C
`define CUBE_LUT_3E2B 16'h3B4D
`define CUBE_LUT_3E2C 16'h3B4D
`define CUBE_LUT_3E2D 16'h3B4D
`define CUBE_LUT_3E2E 16'h3B4E
`define CUBE_LUT_3E2F 16'h3B4E
`define CUBE_LUT_3E30 16'h3B4E
`define CUBE_LUT_3E31 16'h3B4F
`define CUBE_LUT_3E32 16'h3B4F
`define CUBE_LUT_3E33 16'h3B4F
`define CUBE_LUT_3E34 16'h3B50
`define CUBE_LUT_3E35 16'h3B50
`define CUBE_LUT_3E36 16'h3B50
`define CUBE_LUT_3E37 16'h3B51
`define CUBE_LUT_3E38 16'h3B51
`define CUBE_LUT_3E39 16'h3B51
`define CUBE_LUT_3E3A 16'h3B52
`define CUBE_LUT_3E3B 16'h3B52
`define CUBE_LUT_3E3C 16'h3B52
`define CUBE_LUT_3E3D 16'h3B53
`define CUBE_LUT_3E3E 16'h3B53
`define CUBE_LUT_3E3F 16'h3B53
`define CUBE_LUT_3E40 16'h3B54
`define CUBE_LUT_3E41 16'h3B54
`define CUBE_LUT_3E42 16'h3B54
`define CUBE_LUT_3E43 16'h3B55
`define CUBE_LUT_3E44 16'h3B55
`define CUBE_LUT_3E45 16'h3B55
`define CUBE_LUT_3E46 16'h3B56
`define CUBE_LUT_3E47 16'h3B56
`define CUBE_LUT_3E48 16'h3B56
`define CUBE_LUT_3E49 16'h3B56
`define CUBE_LUT_3E4A 16'h3B57
`define CUBE_LUT_3E4B 16'h3B57
`define CUBE_LUT_3E4C 16'h3B57
`define CUBE_LUT_3E4D 16'h3B58
`define CUBE_LUT_3E4E 16'h3B58
`define CUBE_LUT_3E4F 16'h3B58
`define CUBE_LUT_3E50 16'h3B59
`define CUBE_LUT_3E51 16'h3B59
`define CUBE_LUT_3E52 16'h3B59
`define CUBE_LUT_3E53 16'h3B5A
`define CUBE_LUT_3E54 16'h3B5A
`define CUBE_LUT_3E55 16'h3B5A
`define CUBE_LUT_3E56 16'h3B5B
`define CUBE_LUT_3E57 16'h3B5B
`define CUBE_LUT_3E58 16'h3B5B
`define CUBE_LUT_3E59 16'h3B5B
`define CUBE_LUT_3E5A 16'h3B5C
`define CUBE_LUT_3E5B 16'h3B5C
`define CUBE_LUT_3E5C 16'h3B5C
`define CUBE_LUT_3E5D 16'h3B5D
`define CUBE_LUT_3E5E 16'h3B5D
`define CUBE_LUT_3E5F 16'h3B5D
`define CUBE_LUT_3E60 16'h3B5E
`define CUBE_LUT_3E61 16'h3B5E
`define CUBE_LUT_3E62 16'h3B5E
`define CUBE_LUT_3E63 16'h3B5F
`define CUBE_LUT_3E64 16'h3B5F
`define CUBE_LUT_3E65 16'h3B5F
`define CUBE_LUT_3E66 16'h3B5F
`define CUBE_LUT_3E67 16'h3B60
`define CUBE_LUT_3E68 16'h3B60
`define CUBE_LUT_3E69 16'h3B60
`define CUBE_LUT_3E6A 16'h3B61
`define CUBE_LUT_3E6B 16'h3B61
`define CUBE_LUT_3E6C 16'h3B61
`define CUBE_LUT_3E6D 16'h3B62
`define CUBE_LUT_3E6E 16'h3B62
`define CUBE_LUT_3E6F 16'h3B62
`define CUBE_LUT_3E70 16'h3B62
`define CUBE_LUT_3E71 16'h3B63
`define CUBE_LUT_3E72 16'h3B63
`define CUBE_LUT_3E73 16'h3B63
`define CUBE_LUT_3E74 16'h3B64
`define CUBE_LUT_3E75 16'h3B64
`define CUBE_LUT_3E76 16'h3B64
`define CUBE_LUT_3E77 16'h3B65
`define CUBE_LUT_3E78 16'h3B65
`define CUBE_LUT_3E79 16'h3B65
`define CUBE_LUT_3E7A 16'h3B65
`define CUBE_LUT_3E7B 16'h3B66
`define CUBE_LUT_3E7C 16'h3B66
`define CUBE_LUT_3E7D 16'h3B66
`define CUBE_LUT_3E7E 16'h3B67
`define CUBE_LUT_3E7F 16'h3B67
`define CUBE_LUT_3E80 16'h3B67
`define CUBE_LUT_3E81 16'h3B67
`define CUBE_LUT_3E82 16'h3B68
`define CUBE_LUT_3E83 16'h3B68
`define CUBE_LUT_3E84 16'h3B68
`define CUBE_LUT_3E85 16'h3B69
`define CUBE_LUT_3E86 16'h3B69
`define CUBE_LUT_3E87 16'h3B69
`define CUBE_LUT_3E88 16'h3B69
`define CUBE_LUT_3E89 16'h3B6A
`define CUBE_LUT_3E8A 16'h3B6A
`define CUBE_LUT_3E8B 16'h3B6A
`define CUBE_LUT_3E8C 16'h3B6B
`define CUBE_LUT_3E8D 16'h3B6B
`define CUBE_LUT_3E8E 16'h3B6B
`define CUBE_LUT_3E8F 16'h3B6B
`define CUBE_LUT_3E90 16'h3B6C
`define CUBE_LUT_3E91 16'h3B6C
`define CUBE_LUT_3E92 16'h3B6C
`define CUBE_LUT_3E93 16'h3B6C
`define CUBE_LUT_3E94 16'h3B6D
`define CUBE_LUT_3E95 16'h3B6D
`define CUBE_LUT_3E96 16'h3B6D
`define CUBE_LUT_3E97 16'h3B6E
`define CUBE_LUT_3E98 16'h3B6E
`define CUBE_LUT_3E99 16'h3B6E
`define CUBE_LUT_3E9A 16'h3B6E
`define CUBE_LUT_3E9B 16'h3B6F
`define CUBE_LUT_3E9C 16'h3B6F
`define CUBE_LUT_3E9D 16'h3B6F
`define CUBE_LUT_3E9E 16'h3B70
`define CUBE_LUT_3E9F 16'h3B70
`define CUBE_LUT_3EA0 16'h3B70
`define CUBE_LUT_3EA1 16'h3B70
`define CUBE_LUT_3EA2 16'h3B71
`define CUBE_LUT_3EA3 16'h3B71
`define CUBE_LUT_3EA4 16'h3B71
`define CUBE_LUT_3EA5 16'h3B71
`define CUBE_LUT_3EA6 16'h3B72
`define CUBE_LUT_3EA7 16'h3B72
`define CUBE_LUT_3EA8 16'h3B72
`define CUBE_LUT_3EA9 16'h3B72
`define CUBE_LUT_3EAA 16'h3B73
`define CUBE_LUT_3EAB 16'h3B73
`define CUBE_LUT_3EAC 16'h3B73
`define CUBE_LUT_3EAD 16'h3B74
`define CUBE_LUT_3EAE 16'h3B74
`define CUBE_LUT_3EAF 16'h3B74
`define CUBE_LUT_3EB0 16'h3B74
`define CUBE_LUT_3EB1 16'h3B75
`define CUBE_LUT_3EB2 16'h3B75
`define CUBE_LUT_3EB3 16'h3B75
`define CUBE_LUT_3EB4 16'h3B75
`define CUBE_LUT_3EB5 16'h3B76
`define CUBE_LUT_3EB6 16'h3B76
`define CUBE_LUT_3EB7 16'h3B76
`define CUBE_LUT_3EB8 16'h3B76
`define CUBE_LUT_3EB9 16'h3B77
`define CUBE_LUT_3EBA 16'h3B77
`define CUBE_LUT_3EBB 16'h3B77
`define CUBE_LUT_3EBC 16'h3B77
`define CUBE_LUT_3EBD 16'h3B78
`define CUBE_LUT_3EBE 16'h3B78
`define CUBE_LUT_3EBF 16'h3B78
`define CUBE_LUT_3EC0 16'h3B78
`define CUBE_LUT_3EC1 16'h3B79
`define CUBE_LUT_3EC2 16'h3B79
`define CUBE_LUT_3EC3 16'h3B79
`define CUBE_LUT_3EC4 16'h3B79
`define CUBE_LUT_3EC5 16'h3B7A
`define CUBE_LUT_3EC6 16'h3B7A
`define CUBE_LUT_3EC7 16'h3B7A
`define CUBE_LUT_3EC8 16'h3B7B
`define CUBE_LUT_3EC9 16'h3B7B
`define CUBE_LUT_3ECA 16'h3B7B
`define CUBE_LUT_3ECB 16'h3B7B
`define CUBE_LUT_3ECC 16'h3B7C
`define CUBE_LUT_3ECD 16'h3B7C
`define CUBE_LUT_3ECE 16'h3B7C
`define CUBE_LUT_3ECF 16'h3B7C
`define CUBE_LUT_3ED0 16'h3B7D
`define CUBE_LUT_3ED1 16'h3B7D
`define CUBE_LUT_3ED2 16'h3B7D
`define CUBE_LUT_3ED3 16'h3B7D
`define CUBE_LUT_3ED4 16'h3B7E
`define CUBE_LUT_3ED5 16'h3B7E
`define CUBE_LUT_3ED6 16'h3B7E
`define CUBE_LUT_3ED7 16'h3B7E
`define CUBE_LUT_3ED8 16'h3B7E
`define CUBE_LUT_3ED9 16'h3B7F
`define CUBE_LUT_3EDA 16'h3B7F
`define CUBE_LUT_3EDB 16'h3B7F
`define CUBE_LUT_3EDC 16'h3B7F
`define CUBE_LUT_3EDD 16'h3B80
`define CUBE_LUT_3EDE 16'h3B80
`define CUBE_LUT_3EDF 16'h3B80
`define CUBE_LUT_3EE0 16'h3B80
`define CUBE_LUT_3EE1 16'h3B81
`define CUBE_LUT_3EE2 16'h3B81
`define CUBE_LUT_3EE3 16'h3B81
`define CUBE_LUT_3EE4 16'h3B81
`define CUBE_LUT_3EE5 16'h3B82
`define CUBE_LUT_3EE6 16'h3B82
`define CUBE_LUT_3EE7 16'h3B82
`define CUBE_LUT_3EE8 16'h3B82
`define CUBE_LUT_3EE9 16'h3B83
`define CUBE_LUT_3EEA 16'h3B83
`define CUBE_LUT_3EEB 16'h3B83
`define CUBE_LUT_3EEC 16'h3B83
`define CUBE_LUT_3EED 16'h3B84
`define CUBE_LUT_3EEE 16'h3B84
`define CUBE_LUT_3EEF 16'h3B84
`define CUBE_LUT_3EF0 16'h3B84
`define CUBE_LUT_3EF1 16'h3B84
`define CUBE_LUT_3EF2 16'h3B85
`define CUBE_LUT_3EF3 16'h3B85
`define CUBE_LUT_3EF4 16'h3B85
`define CUBE_LUT_3EF5 16'h3B85
`define CUBE_LUT_3EF6 16'h3B86
`define CUBE_LUT_3EF7 16'h3B86
`define CUBE_LUT_3EF8 16'h3B86
`define CUBE_LUT_3EF9 16'h3B86
`define CUBE_LUT_3EFA 16'h3B87
`define CUBE_LUT_3EFB 16'h3B87
`define CUBE_LUT_3EFC 16'h3B87
`define CUBE_LUT_3EFD 16'h3B87
`define CUBE_LUT_3EFE 16'h3B87
`define CUBE_LUT_3EFF 16'h3B88
`define CUBE_LUT_3F00 16'h3B88
`define CUBE_LUT_3F01 16'h3B88
`define CUBE_LUT_3F02 16'h3B88
`define CUBE_LUT_3F03 16'h3B89
`define CUBE_LUT_3F04 16'h3B89
`define CUBE_LUT_3F05 16'h3B89
`define CUBE_LUT_3F06 16'h3B89
`define CUBE_LUT_3F07 16'h3B8A
`define CUBE_LUT_3F08 16'h3B8A
`define CUBE_LUT_3F09 16'h3B8A
`define CUBE_LUT_3F0A 16'h3B8A
`define CUBE_LUT_3F0B 16'h3B8A
`define CUBE_LUT_3F0C 16'h3B8B
`define CUBE_LUT_3F0D 16'h3B8B
`define CUBE_LUT_3F0E 16'h3B8B
`define CUBE_LUT_3F0F 16'h3B8B
`define CUBE_LUT_3F10 16'h3B8C
`define CUBE_LUT_3F11 16'h3B8C
`define CUBE_LUT_3F12 16'h3B8C
`define CUBE_LUT_3F13 16'h3B8C
`define CUBE_LUT_3F14 16'h3B8C
`define CUBE_LUT_3F15 16'h3B8D
`define CUBE_LUT_3F16 16'h3B8D
`define CUBE_LUT_3F17 16'h3B8D
`define CUBE_LUT_3F18 16'h3B8D
`define CUBE_LUT_3F19 16'h3B8D
`define CUBE_LUT_3F1A 16'h3B8E
`define CUBE_LUT_3F1B 16'h3B8E
`define CUBE_LUT_3F1C 16'h3B8E
`define CUBE_LUT_3F1D 16'h3B8E
`define CUBE_LUT_3F1E 16'h3B8F
`define CUBE_LUT_3F1F 16'h3B8F
`define CUBE_LUT_3F20 16'h3B8F
`define CUBE_LUT_3F21 16'h3B8F
`define CUBE_LUT_3F22 16'h3B8F
`define CUBE_LUT_3F23 16'h3B90
`define CUBE_LUT_3F24 16'h3B90
`define CUBE_LUT_3F25 16'h3B90
`define CUBE_LUT_3F26 16'h3B90
`define CUBE_LUT_3F27 16'h3B91
`define CUBE_LUT_3F28 16'h3B91
`define CUBE_LUT_3F29 16'h3B91
`define CUBE_LUT_3F2A 16'h3B91
`define CUBE_LUT_3F2B 16'h3B91
`define CUBE_LUT_3F2C 16'h3B92
`define CUBE_LUT_3F2D 16'h3B92
`define CUBE_LUT_3F2E 16'h3B92
`define CUBE_LUT_3F2F 16'h3B92
`define CUBE_LUT_3F30 16'h3B92
`define CUBE_LUT_3F31 16'h3B93
`define CUBE_LUT_3F32 16'h3B93
`define CUBE_LUT_3F33 16'h3B93
`define CUBE_LUT_3F34 16'h3B93
`define CUBE_LUT_3F35 16'h3B93
`define CUBE_LUT_3F36 16'h3B94
`define CUBE_LUT_3F37 16'h3B94
`define CUBE_LUT_3F38 16'h3B94
`define CUBE_LUT_3F39 16'h3B94
`define CUBE_LUT_3F3A 16'h3B94
`define CUBE_LUT_3F3B 16'h3B95
`define CUBE_LUT_3F3C 16'h3B95
`define CUBE_LUT_3F3D 16'h3B95
`define CUBE_LUT_3F3E 16'h3B95
`define CUBE_LUT_3F3F 16'h3B95
`define CUBE_LUT_3F40 16'h3B96
`define CUBE_LUT_3F41 16'h3B96
`define CUBE_LUT_3F42 16'h3B96
`define CUBE_LUT_3F43 16'h3B96
`define CUBE_LUT_3F44 16'h3B96
`define CUBE_LUT_3F45 16'h3B97
`define CUBE_LUT_3F46 16'h3B97
`define CUBE_LUT_3F47 16'h3B97
`define CUBE_LUT_3F48 16'h3B97
`define CUBE_LUT_3F49 16'h3B97
`define CUBE_LUT_3F4A 16'h3B98
`define CUBE_LUT_3F4B 16'h3B98
`define CUBE_LUT_3F4C 16'h3B98
`define CUBE_LUT_3F4D 16'h3B98
`define CUBE_LUT_3F4E 16'h3B98
`define CUBE_LUT_3F4F 16'h3B99
`define CUBE_LUT_3F50 16'h3B99
`define CUBE_LUT_3F51 16'h3B99
`define CUBE_LUT_3F52 16'h3B99
`define CUBE_LUT_3F53 16'h3B99
`define CUBE_LUT_3F54 16'h3B9A
`define CUBE_LUT_3F55 16'h3B9A
`define CUBE_LUT_3F56 16'h3B9A
`define CUBE_LUT_3F57 16'h3B9A
`define CUBE_LUT_3F58 16'h3B9A
`define CUBE_LUT_3F59 16'h3B9B
`define CUBE_LUT_3F5A 16'h3B9B
`define CUBE_LUT_3F5B 16'h3B9B
`define CUBE_LUT_3F5C 16'h3B9B
`define CUBE_LUT_3F5D 16'h3B9B
`define CUBE_LUT_3F5E 16'h3B9C
`define CUBE_LUT_3F5F 16'h3B9C
`define CUBE_LUT_3F60 16'h3B9C
`define CUBE_LUT_3F61 16'h3B9C
`define CUBE_LUT_3F62 16'h3B9C
`define CUBE_LUT_3F63 16'h3B9D
`define CUBE_LUT_3F64 16'h3B9D
`define CUBE_LUT_3F65 16'h3B9D
`define CUBE_LUT_3F66 16'h3B9D
`define CUBE_LUT_3F67 16'h3B9D
`define CUBE_LUT_3F68 16'h3B9D
`define CUBE_LUT_3F69 16'h3B9E
`define CUBE_LUT_3F6A 16'h3B9E
`define CUBE_LUT_3F6B 16'h3B9E
`define CUBE_LUT_3F6C 16'h3B9E
`define CUBE_LUT_3F6D 16'h3B9E
`define CUBE_LUT_3F6E 16'h3B9F
`define CUBE_LUT_3F6F 16'h3B9F
`define CUBE_LUT_3F70 16'h3B9F
`define CUBE_LUT_3F71 16'h3B9F
`define CUBE_LUT_3F72 16'h3B9F
`define CUBE_LUT_3F73 16'h3BA0
`define CUBE_LUT_3F74 16'h3BA0
`define CUBE_LUT_3F75 16'h3BA0
`define CUBE_LUT_3F76 16'h3BA0
`define CUBE_LUT_3F77 16'h3BA0
`define CUBE_LUT_3F78 16'h3BA0
`define CUBE_LUT_3F79 16'h3BA1
`define CUBE_LUT_3F7A 16'h3BA1
`define CUBE_LUT_3F7B 16'h3BA1
`define CUBE_LUT_3F7C 16'h3BA1
`define CUBE_LUT_3F7D 16'h3BA1
`define CUBE_LUT_3F7E 16'h3BA2
`define CUBE_LUT_3F7F 16'h3BA2
`define CUBE_LUT_3F80 16'h3BA2
`define CUBE_LUT_3F81 16'h3BA2
`define CUBE_LUT_3F82 16'h3BA2
`define CUBE_LUT_3F83 16'h3BA2
`define CUBE_LUT_3F84 16'h3BA3
`define CUBE_LUT_3F85 16'h3BA3
`define CUBE_LUT_3F86 16'h3BA3
`define CUBE_LUT_3F87 16'h3BA3
`define CUBE_LUT_3F88 16'h3BA3
`define CUBE_LUT_3F89 16'h3BA3
`define CUBE_LUT_3F8A 16'h3BA4
`define CUBE_LUT_3F8B 16'h3BA4
`define CUBE_LUT_3F8C 16'h3BA4
`define CUBE_LUT_3F8D 16'h3BA4
`define CUBE_LUT_3F8E 16'h3BA4
`define CUBE_LUT_3F8F 16'h3BA5
`define CUBE_LUT_3F90 16'h3BA5
`define CUBE_LUT_3F91 16'h3BA5
`define CUBE_LUT_3F92 16'h3BA5
`define CUBE_LUT_3F93 16'h3BA5
`define CUBE_LUT_3F94 16'h3BA5
`define CUBE_LUT_3F95 16'h3BA6
`define CUBE_LUT_3F96 16'h3BA6
`define CUBE_LUT_3F97 16'h3BA6
`define CUBE_LUT_3F98 16'h3BA6
`define CUBE_LUT_3F99 16'h3BA6
`define CUBE_LUT_3F9A 16'h3BA6
`define CUBE_LUT_3F9B 16'h3BA7
`define CUBE_LUT_3F9C 16'h3BA7
`define CUBE_LUT_3F9D 16'h3BA7
`define CUBE_LUT_3F9E 16'h3BA7
`define CUBE_LUT_3F9F 16'h3BA7
`define CUBE_LUT_3FA0 16'h3BA7
`define CUBE_LUT_3FA1 16'h3BA8
`define CUBE_LUT_3FA2 16'h3BA8
`define CUBE_LUT_3FA3 16'h3BA8
`define CUBE_LUT_3FA4 16'h3BA8
`define CUBE_LUT_3FA5 16'h3BA8
`define CUBE_LUT_3FA6 16'h3BA8
`define CUBE_LUT_3FA7 16'h3BA9
`define CUBE_LUT_3FA8 16'h3BA9
`define CUBE_LUT_3FA9 16'h3BA9
`define CUBE_LUT_3FAA 16'h3BA9
`define CUBE_LUT_3FAB 16'h3BA9
`define CUBE_LUT_3FAC 16'h3BA9
`define CUBE_LUT_3FAD 16'h3BAA
`define CUBE_LUT_3FAE 16'h3BAA
`define CUBE_LUT_3FAF 16'h3BAA
`define CUBE_LUT_3FB0 16'h3BAA
`define CUBE_LUT_3FB1 16'h3BAA
`define CUBE_LUT_3FB2 16'h3BAA
`define CUBE_LUT_3FB3 16'h3BAB
`define CUBE_LUT_3FB4 16'h3BAB
`define CUBE_LUT_3FB5 16'h3BAB
`define CUBE_LUT_3FB6 16'h3BAB
`define CUBE_LUT_3FB7 16'h3BAB
`define CUBE_LUT_3FB8 16'h3BAB
`define CUBE_LUT_3FB9 16'h3BAC
`define CUBE_LUT_3FBA 16'h3BAC
`define CUBE_LUT_3FBB 16'h3BAC
`define CUBE_LUT_3FBC 16'h3BAC
`define CUBE_LUT_3FBD 16'h3BAC
`define CUBE_LUT_3FBE 16'h3BAC
`define CUBE_LUT_3FBF 16'h3BAD
`define CUBE_LUT_3FC0 16'h3BAD
`define CUBE_LUT_3FC1 16'h3BAD
`define CUBE_LUT_3FC2 16'h3BAD
`define CUBE_LUT_3FC3 16'h3BAD
`define CUBE_LUT_3FC4 16'h3BAD
`define CUBE_LUT_3FC5 16'h3BAE
`define CUBE_LUT_3FC6 16'h3BAE
`define CUBE_LUT_3FC7 16'h3BAE
`define CUBE_LUT_3FC8 16'h3BAE
`define CUBE_LUT_3FC9 16'h3BAE
`define CUBE_LUT_3FCA 16'h3BAE
`define CUBE_LUT_3FCB 16'h3BAE
`define CUBE_LUT_3FCC 16'h3BAF
`define CUBE_LUT_3FCD 16'h3BAF
`define CUBE_LUT_3FCE 16'h3BAF
`define CUBE_LUT_3FCF 16'h3BAF
`define CUBE_LUT_3FD0 16'h3BAF
`define CUBE_LUT_3FD1 16'h3BAF
`define CUBE_LUT_3FD2 16'h3BB0
`define CUBE_LUT_3FD3 16'h3BB0
`define CUBE_LUT_3FD4 16'h3BB0
`define CUBE_LUT_3FD5 16'h3BB0
`define CUBE_LUT_3FD6 16'h3BB0
`define CUBE_LUT_3FD7 16'h3BB0
`define CUBE_LUT_3FD8 16'h3BB0
`define CUBE_LUT_3FD9 16'h3BB1
`define CUBE_LUT_3FDA 16'h3BB1
`define CUBE_LUT_3FDB 16'h3BB1
`define CUBE_LUT_3FDC 16'h3BB1
`define CUBE_LUT_3FDD 16'h3BB1
`define CUBE_LUT_3FDE 16'h3BB1
`define CUBE_LUT_3FDF 16'h3BB2
`define CUBE_LUT_3FE0 16'h3BB2
`define CUBE_LUT_3FE1 16'h3BB2
`define CUBE_LUT_3FE2 16'h3BB2
`define CUBE_LUT_3FE3 16'h3BB2
`define CUBE_LUT_3FE4 16'h3BB2
`define CUBE_LUT_3FE5 16'h3BB2
`define CUBE_LUT_3FE6 16'h3BB3
`define CUBE_LUT_3FE7 16'h3BB3
`define CUBE_LUT_3FE8 16'h3BB3
`define CUBE_LUT_3FE9 16'h3BB3
`define CUBE_LUT_3FEA 16'h3BB3
`define CUBE_LUT_3FEB 16'h3BB3
`define CUBE_LUT_3FEC 16'h3BB3
`define CUBE_LUT_3FED 16'h3BB4
`define CUBE_LUT_3FEE 16'h3BB4
`define CUBE_LUT_3FEF 16'h3BB4
`define CUBE_LUT_3FF0 16'h3BB4
`define CUBE_LUT_3FF1 16'h3BB4
`define CUBE_LUT_3FF2 16'h3BB4
`define CUBE_LUT_3FF3 16'h3BB4
`define CUBE_LUT_3FF4 16'h3BB5
`define CUBE_LUT_3FF5 16'h3BB5
`define CUBE_LUT_3FF6 16'h3BB5
`define CUBE_LUT_3FF7 16'h3BB5
`define CUBE_LUT_3FF8 16'h3BB5
`define CUBE_LUT_3FF9 16'h3BB5
`define CUBE_LUT_3FFA 16'h3BB5
`define CUBE_LUT_3FFB 16'h3BB6
`define CUBE_LUT_3FFC 16'h3BB6
`define CUBE_LUT_3FFD 16'h3BB6
`define CUBE_LUT_3FFE 16'h3BB6
`define CUBE_LUT_3FFF 16'h3BB6
`define CUBE_LUT_4000 16'h3BB6
`define CUBE_LUT_4001 16'h3BB7
`define CUBE_LUT_4002 16'h3BB7
`define CUBE_LUT_4003 16'h3BB7
`define CUBE_LUT_4004 16'h3BB7
`define CUBE_LUT_4005 16'h3BB8
`define CUBE_LUT_4006 16'h3BB8
`define CUBE_LUT_4007 16'h3BB8
`define CUBE_LUT_4008 16'h3BB9
`define CUBE_LUT_4009 16'h3BB9
`define CUBE_LUT_400A 16'h3BB9
`define CUBE_LUT_400B 16'h3BB9
`define CUBE_LUT_400C 16'h3BBA
`define CUBE_LUT_400D 16'h3BBA
`define CUBE_LUT_400E 16'h3BBA
`define CUBE_LUT_400F 16'h3BBA
`define CUBE_LUT_4010 16'h3BBB
`define CUBE_LUT_4011 16'h3BBB
`define CUBE_LUT_4012 16'h3BBB
`define CUBE_LUT_4013 16'h3BBC
`define CUBE_LUT_4014 16'h3BBC
`define CUBE_LUT_4015 16'h3BBC
`define CUBE_LUT_4016 16'h3BBC
`define CUBE_LUT_4017 16'h3BBD
`define CUBE_LUT_4018 16'h3BBD
`define CUBE_LUT_4019 16'h3BBD
`define CUBE_LUT_401A 16'h3BBD
`define CUBE_LUT_401B 16'h3BBE
`define CUBE_LUT_401C 16'h3BBE
`define CUBE_LUT_401D 16'h3BBE
`define CUBE_LUT_401E 16'h3BBE
`define CUBE_LUT_401F 16'h3BBF
`define CUBE_LUT_4020 16'h3BBF
`define CUBE_LUT_4021 16'h3BBF
`define CUBE_LUT_4022 16'h3BBF
`define CUBE_LUT_4023 16'h3BC0
`define CUBE_LUT_4024 16'h3BC0
`define CUBE_LUT_4025 16'h3BC0
`define CUBE_LUT_4026 16'h3BC0
`define CUBE_LUT_4027 16'h3BC1
`define CUBE_LUT_4028 16'h3BC1
`define CUBE_LUT_4029 16'h3BC1
`define CUBE_LUT_402A 16'h3BC1
`define CUBE_LUT_402B 16'h3BC2
`define CUBE_LUT_402C 16'h3BC2
`define CUBE_LUT_402D 16'h3BC2
`define CUBE_LUT_402E 16'h3BC2
`define CUBE_LUT_402F 16'h3BC2
`define CUBE_LUT_4030 16'h3BC3
`define CUBE_LUT_4031 16'h3BC3
`define CUBE_LUT_4032 16'h3BC3
`define CUBE_LUT_4033 16'h3BC3
`define CUBE_LUT_4034 16'h3BC4
`define CUBE_LUT_4035 16'h3BC4
`define CUBE_LUT_4036 16'h3BC4
`define CUBE_LUT_4037 16'h3BC4
`define CUBE_LUT_4038 16'h3BC5
`define CUBE_LUT_4039 16'h3BC5
`define CUBE_LUT_403A 16'h3BC5
`define CUBE_LUT_403B 16'h3BC5
`define CUBE_LUT_403C 16'h3BC6
`define CUBE_LUT_403D 16'h3BC6
`define CUBE_LUT_403E 16'h3BC6
`define CUBE_LUT_403F 16'h3BC6
`define CUBE_LUT_4040 16'h3BC6
`define CUBE_LUT_4041 16'h3BC7
`define CUBE_LUT_4042 16'h3BC7
`define CUBE_LUT_4043 16'h3BC7
`define CUBE_LUT_4044 16'h3BC7
`define CUBE_LUT_4045 16'h3BC7
`define CUBE_LUT_4046 16'h3BC8
`define CUBE_LUT_4047 16'h3BC8
`define CUBE_LUT_4048 16'h3BC8
`define CUBE_LUT_4049 16'h3BC8
`define CUBE_LUT_404A 16'h3BC9
`define CUBE_LUT_404B 16'h3BC9
`define CUBE_LUT_404C 16'h3BC9
`define CUBE_LUT_404D 16'h3BC9
`define CUBE_LUT_404E 16'h3BC9
`define CUBE_LUT_404F 16'h3BCA
`define CUBE_LUT_4050 16'h3BCA
`define CUBE_LUT_4051 16'h3BCA
`define CUBE_LUT_4052 16'h3BCA
`define CUBE_LUT_4053 16'h3BCA
`define CUBE_LUT_4054 16'h3BCB
`define CUBE_LUT_4055 16'h3BCB
`define CUBE_LUT_4056 16'h3BCB
`define CUBE_LUT_4057 16'h3BCB
`define CUBE_LUT_4058 16'h3BCB
`define CUBE_LUT_4059 16'h3BCC
`define CUBE_LUT_405A 16'h3BCC
`define CUBE_LUT_405B 16'h3BCC
`define CUBE_LUT_405C 16'h3BCC
`define CUBE_LUT_405D 16'h3BCC
`define CUBE_LUT_405E 16'h3BCD
`define CUBE_LUT_405F 16'h3BCD
`define CUBE_LUT_4060 16'h3BCD
`define CUBE_LUT_4061 16'h3BCD
`define CUBE_LUT_4062 16'h3BCD
`define CUBE_LUT_4063 16'h3BCE
`define CUBE_LUT_4064 16'h3BCE
`define CUBE_LUT_4065 16'h3BCE
`define CUBE_LUT_4066 16'h3BCE
`define CUBE_LUT_4067 16'h3BCE
`define CUBE_LUT_4068 16'h3BCF
`define CUBE_LUT_4069 16'h3BCF
`define CUBE_LUT_406A 16'h3BCF
`define CUBE_LUT_406B 16'h3BCF
`define CUBE_LUT_406C 16'h3BCF
`define CUBE_LUT_406D 16'h3BD0
`define CUBE_LUT_406E 16'h3BD0
`define CUBE_LUT_406F 16'h3BD0
`define CUBE_LUT_4070 16'h3BD0
`define CUBE_LUT_4071 16'h3BD0
`define CUBE_LUT_4072 16'h3BD0
`define CUBE_LUT_4073 16'h3BD1
`define CUBE_LUT_4074 16'h3BD1
`define CUBE_LUT_4075 16'h3BD1
`define CUBE_LUT_4076 16'h3BD1
`define CUBE_LUT_4077 16'h3BD1
`define CUBE_LUT_4078 16'h3BD2
`define CUBE_LUT_4079 16'h3BD2
`define CUBE_LUT_407A 16'h3BD2
`define CUBE_LUT_407B 16'h3BD2
`define CUBE_LUT_407C 16'h3BD2
`define CUBE_LUT_407D 16'h3BD2
`define CUBE_LUT_407E 16'h3BD3
`define CUBE_LUT_407F 16'h3BD3
`define CUBE_LUT_4080 16'h3BD3
`define CUBE_LUT_4081 16'h3BD3
`define CUBE_LUT_4082 16'h3BD3
`define CUBE_LUT_4083 16'h3BD4
`define CUBE_LUT_4084 16'h3BD4
`define CUBE_LUT_4085 16'h3BD4
`define CUBE_LUT_4086 16'h3BD4
`define CUBE_LUT_4087 16'h3BD4
`define CUBE_LUT_4088 16'h3BD4
`define CUBE_LUT_4089 16'h3BD5
`define CUBE_LUT_408A 16'h3BD5
`define CUBE_LUT_408B 16'h3BD5
`define CUBE_LUT_408C 16'h3BD5
`define CUBE_LUT_408D 16'h3BD5
`define CUBE_LUT_408E 16'h3BD5
`define CUBE_LUT_408F 16'h3BD6
`define CUBE_LUT_4090 16'h3BD6
`define CUBE_LUT_4091 16'h3BD6
`define CUBE_LUT_4092 16'h3BD6
`define CUBE_LUT_4093 16'h3BD6
`define CUBE_LUT_4094 16'h3BD6
`define CUBE_LUT_4095 16'h3BD7
`define CUBE_LUT_4096 16'h3BD7
`define CUBE_LUT_4097 16'h3BD7
`define CUBE_LUT_4098 16'h3BD7
`define CUBE_LUT_4099 16'h3BD7
`define CUBE_LUT_409A 16'h3BD7
`define CUBE_LUT_409B 16'h3BD7
`define CUBE_LUT_409C 16'h3BD8
`define CUBE_LUT_409D 16'h3BD8
`define CUBE_LUT_409E 16'h3BD8
`define CUBE_LUT_409F 16'h3BD8
`define CUBE_LUT_40A0 16'h3BD8
`define CUBE_LUT_40A1 16'h3BD8
`define CUBE_LUT_40A2 16'h3BD9
`define CUBE_LUT_40A3 16'h3BD9
`define CUBE_LUT_40A4 16'h3BD9
`define CUBE_LUT_40A5 16'h3BD9
`define CUBE_LUT_40A6 16'h3BD9
`define CUBE_LUT_40A7 16'h3BD9
`define CUBE_LUT_40A8 16'h3BD9
`define CUBE_LUT_40A9 16'h3BDA
`define CUBE_LUT_40AA 16'h3BDA
`define CUBE_LUT_40AB 16'h3BDA
`define CUBE_LUT_40AC 16'h3BDA
`define CUBE_LUT_40AD 16'h3BDA
`define CUBE_LUT_40AE 16'h3BDA
`define CUBE_LUT_40AF 16'h3BDA
`define CUBE_LUT_40B0 16'h3BDB
`define CUBE_LUT_40B1 16'h3BDB
`define CUBE_LUT_40B2 16'h3BDB
`define CUBE_LUT_40B3 16'h3BDB
`define CUBE_LUT_40B4 16'h3BDB
`define CUBE_LUT_40B5 16'h3BDB
`define CUBE_LUT_40B6 16'h3BDB
`define CUBE_LUT_40B7 16'h3BDC
`define CUBE_LUT_40B8 16'h3BDC
`define CUBE_LUT_40B9 16'h3BDC
`define CUBE_LUT_40BA 16'h3BDC
`define CUBE_LUT_40BB 16'h3BDC
`define CUBE_LUT_40BC 16'h3BDC
`define CUBE_LUT_40BD 16'h3BDC
`define CUBE_LUT_40BE 16'h3BDD
`define CUBE_LUT_40BF 16'h3BDD
`define CUBE_LUT_40C0 16'h3BDD
`define CUBE_LUT_40C1 16'h3BDD
`define CUBE_LUT_40C2 16'h3BDD
`define CUBE_LUT_40C3 16'h3BDD
`define CUBE_LUT_40C4 16'h3BDD
`define CUBE_LUT_40C5 16'h3BDE
`define CUBE_LUT_40C6 16'h3BDE
`define CUBE_LUT_40C7 16'h3BDE
`define CUBE_LUT_40C8 16'h3BDE
`define CUBE_LUT_40C9 16'h3BDE
`define CUBE_LUT_40CA 16'h3BDE
`define CUBE_LUT_40CB 16'h3BDE
`define CUBE_LUT_40CC 16'h3BDE
`define CUBE_LUT_40CD 16'h3BDF
`define CUBE_LUT_40CE 16'h3BDF
`define CUBE_LUT_40CF 16'h3BDF
`define CUBE_LUT_40D0 16'h3BDF
`define CUBE_LUT_40D1 16'h3BDF
`define CUBE_LUT_40D2 16'h3BDF
`define CUBE_LUT_40D3 16'h3BDF
`define CUBE_LUT_40D4 16'h3BDF
`define CUBE_LUT_40D5 16'h3BE0
`define CUBE_LUT_40D6 16'h3BE0
`define CUBE_LUT_40D7 16'h3BE0
`define CUBE_LUT_40D8 16'h3BE0
`define CUBE_LUT_40D9 16'h3BE0
`define CUBE_LUT_40DA 16'h3BE0
`define CUBE_LUT_40DB 16'h3BE0
`define CUBE_LUT_40DC 16'h3BE0
`define CUBE_LUT_40DD 16'h3BE1
`define CUBE_LUT_40DE 16'h3BE1
`define CUBE_LUT_40DF 16'h3BE1
`define CUBE_LUT_40E0 16'h3BE1
`define CUBE_LUT_40E1 16'h3BE1
`define CUBE_LUT_40E2 16'h3BE1
`define CUBE_LUT_40E3 16'h3BE1
`define CUBE_LUT_40E4 16'h3BE1
`define CUBE_LUT_40E5 16'h3BE2
`define CUBE_LUT_40E6 16'h3BE2
`define CUBE_LUT_40E7 16'h3BE2
`define CUBE_LUT_40E8 16'h3BE2
`define CUBE_LUT_40E9 16'h3BE2
`define CUBE_LUT_40EA 16'h3BE2
`define CUBE_LUT_40EB 16'h3BE2
`define CUBE_LUT_40EC 16'h3BE2
`define CUBE_LUT_40ED 16'h3BE2
`define CUBE_LUT_40EE 16'h3BE3
`define CUBE_LUT_40EF 16'h3BE3
`define CUBE_LUT_40F0 16'h3BE3
`define CUBE_LUT_40F1 16'h3BE3
`define CUBE_LUT_40F2 16'h3BE3
`define CUBE_LUT_40F3 16'h3BE3
`define CUBE_LUT_40F4 16'h3BE3
`define CUBE_LUT_40F5 16'h3BE3
`define CUBE_LUT_40F6 16'h3BE4
`define CUBE_LUT_40F7 16'h3BE4
`define CUBE_LUT_40F8 16'h3BE4
`define CUBE_LUT_40F9 16'h3BE4
`define CUBE_LUT_40FA 16'h3BE4
`define CUBE_LUT_40FB 16'h3BE4
`define CUBE_LUT_40FC 16'h3BE4
`define CUBE_LUT_40FD 16'h3BE4
`define CUBE_LUT_40FE 16'h3BE4
`define CUBE_LUT_40FF 16'h3BE4
`define CUBE_LUT_4100 16'h3BE5
`define CUBE_LUT_4101 16'h3BE5
`define CUBE_LUT_4102 16'h3BE5
`define CUBE_LUT_4103 16'h3BE5
`define CUBE_LUT_4104 16'h3BE5
`define CUBE_LUT_4105 16'h3BE5
`define CUBE_LUT_4106 16'h3BE5
`define CUBE_LUT_4107 16'h3BE5
`define CUBE_LUT_4108 16'h3BE5
`define CUBE_LUT_4109 16'h3BE6
`define CUBE_LUT_410A 16'h3BE6
`define CUBE_LUT_410B 16'h3BE6
`define CUBE_LUT_410C 16'h3BE6
`define CUBE_LUT_410D 16'h3BE6
`define CUBE_LUT_410E 16'h3BE6
`define CUBE_LUT_410F 16'h3BE6
`define CUBE_LUT_4110 16'h3BE6
`define CUBE_LUT_4111 16'h3BE6
`define CUBE_LUT_4112 16'h3BE6
`define CUBE_LUT_4113 16'h3BE7
`define CUBE_LUT_4114 16'h3BE7
`define CUBE_LUT_4115 16'h3BE7
`define CUBE_LUT_4116 16'h3BE7
`define CUBE_LUT_4117 16'h3BE7
`define CUBE_LUT_4118 16'h3BE7
`define CUBE_LUT_4119 16'h3BE7
`define CUBE_LUT_411A 16'h3BE7
`define CUBE_LUT_411B 16'h3BE7
`define CUBE_LUT_411C 16'h3BE7
`define CUBE_LUT_411D 16'h3BE8
`define CUBE_LUT_411E 16'h3BE8
`define CUBE_LUT_411F 16'h3BE8
`define CUBE_LUT_4120 16'h3BE8
`define CUBE_LUT_4121 16'h3BE8
`define CUBE_LUT_4122 16'h3BE8
`define CUBE_LUT_4123 16'h3BE8
`define CUBE_LUT_4124 16'h3BE8
`define CUBE_LUT_4125 16'h3BE8
`define CUBE_LUT_4126 16'h3BE8
`define CUBE_LUT_4127 16'h3BE8
`define CUBE_LUT_4128 16'h3BE9
`define CUBE_LUT_4129 16'h3BE9
`define CUBE_LUT_412A 16'h3BE9
`define CUBE_LUT_412B 16'h3BE9
`define CUBE_LUT_412C 16'h3BE9
`define CUBE_LUT_412D 16'h3BE9
`define CUBE_LUT_412E 16'h3BE9
`define CUBE_LUT_412F 16'h3BE9
`define CUBE_LUT_4130 16'h3BE9
`define CUBE_LUT_4131 16'h3BE9
`define CUBE_LUT_4132 16'h3BE9
`define CUBE_LUT_4133 16'h3BEA
`define CUBE_LUT_4134 16'h3BEA
`define CUBE_LUT_4135 16'h3BEA
`define CUBE_LUT_4136 16'h3BEA
`define CUBE_LUT_4137 16'h3BEA
`define CUBE_LUT_4138 16'h3BEA
`define CUBE_LUT_4139 16'h3BEA
`define CUBE_LUT_413A 16'h3BEA
`define CUBE_LUT_413B 16'h3BEA
`define CUBE_LUT_413C 16'h3BEA
`define CUBE_LUT_413D 16'h3BEA
`define CUBE_LUT_413E 16'h3BEA
`define CUBE_LUT_413F 16'h3BEB
`define CUBE_LUT_4140 16'h3BEB
`define CUBE_LUT_4141 16'h3BEB
`define CUBE_LUT_4142 16'h3BEB
`define CUBE_LUT_4143 16'h3BEB
`define CUBE_LUT_4144 16'h3BEB
`define CUBE_LUT_4145 16'h3BEB
`define CUBE_LUT_4146 16'h3BEB
`define CUBE_LUT_4147 16'h3BEB
`define CUBE_LUT_4148 16'h3BEB
`define CUBE_LUT_4149 16'h3BEB
`define CUBE_LUT_414A 16'h3BEB
`define CUBE_LUT_414B 16'h3BEC
`define CUBE_LUT_414C 16'h3BEC
`define CUBE_LUT_414D 16'h3BEC
`define CUBE_LUT_414E 16'h3BEC
`define CUBE_LUT_414F 16'h3BEC
`define CUBE_LUT_4150 16'h3BEC
`define CUBE_LUT_4151 16'h3BEC
`define CUBE_LUT_4152 16'h3BEC
`define CUBE_LUT_4153 16'h3BEC
`define CUBE_LUT_4154 16'h3BEC
`define CUBE_LUT_4155 16'h3BEC
`define CUBE_LUT_4156 16'h3BEC
`define CUBE_LUT_4157 16'h3BEC
`define CUBE_LUT_4158 16'h3BED
`define CUBE_LUT_4159 16'h3BED
`define CUBE_LUT_415A 16'h3BED
`define CUBE_LUT_415B 16'h3BED
`define CUBE_LUT_415C 16'h3BED
`define CUBE_LUT_415D 16'h3BED
`define CUBE_LUT_415E 16'h3BED
`define CUBE_LUT_415F 16'h3BED
`define CUBE_LUT_4160 16'h3BED
`define CUBE_LUT_4161 16'h3BED
`define CUBE_LUT_4162 16'h3BED
`define CUBE_LUT_4163 16'h3BED
`define CUBE_LUT_4164 16'h3BED
`define CUBE_LUT_4165 16'h3BED
`define CUBE_LUT_4166 16'h3BEE
`define CUBE_LUT_4167 16'h3BEE
`define CUBE_LUT_4168 16'h3BEE
`define CUBE_LUT_4169 16'h3BEE
`define CUBE_LUT_416A 16'h3BEE
`define CUBE_LUT_416B 16'h3BEE
`define CUBE_LUT_416C 16'h3BEE
`define CUBE_LUT_416D 16'h3BEE
`define CUBE_LUT_416E 16'h3BEE
`define CUBE_LUT_416F 16'h3BEE
`define CUBE_LUT_4170 16'h3BEE
`define CUBE_LUT_4171 16'h3BEE
`define CUBE_LUT_4172 16'h3BEE
`define CUBE_LUT_4173 16'h3BEE
`define CUBE_LUT_4174 16'h3BEF
`define CUBE_LUT_4175 16'h3BEF
`define CUBE_LUT_4176 16'h3BEF
`define CUBE_LUT_4177 16'h3BEF
`define CUBE_LUT_4178 16'h3BEF
`define CUBE_LUT_4179 16'h3BEF
`define CUBE_LUT_417A 16'h3BEF
`define CUBE_LUT_417B 16'h3BEF
`define CUBE_LUT_417C 16'h3BEF
`define CUBE_LUT_417D 16'h3BEF
`define CUBE_LUT_417E 16'h3BEF
`define CUBE_LUT_417F 16'h3BEF
`define CUBE_LUT_4180 16'h3BEF
`define CUBE_LUT_4181 16'h3BEF
`define CUBE_LUT_4182 16'h3BEF
`define CUBE_LUT_4183 16'h3BF0
`define CUBE_LUT_4184 16'h3BF0
`define CUBE_LUT_4185 16'h3BF0
`define CUBE_LUT_4186 16'h3BF0
`define CUBE_LUT_4187 16'h3BF0
`define CUBE_LUT_4188 16'h3BF0
`define CUBE_LUT_4189 16'h3BF0
`define CUBE_LUT_418A 16'h3BF0
`define CUBE_LUT_418B 16'h3BF0
`define CUBE_LUT_418C 16'h3BF0
`define CUBE_LUT_418D 16'h3BF0
`define CUBE_LUT_418E 16'h3BF0
`define CUBE_LUT_418F 16'h3BF0
`define CUBE_LUT_4190 16'h3BF0
`define CUBE_LUT_4191 16'h3BF0
`define CUBE_LUT_4192 16'h3BF0
`define CUBE_LUT_4193 16'h3BF1
`define CUBE_LUT_4194 16'h3BF1
`define CUBE_LUT_4195 16'h3BF1
`define CUBE_LUT_4196 16'h3BF1
`define CUBE_LUT_4197 16'h3BF1
`define CUBE_LUT_4198 16'h3BF1
`define CUBE_LUT_4199 16'h3BF1
`define CUBE_LUT_419A 16'h3BF1
`define CUBE_LUT_419B 16'h3BF1
`define CUBE_LUT_419C 16'h3BF1
`define CUBE_LUT_419D 16'h3BF1
`define CUBE_LUT_419E 16'h3BF1
`define CUBE_LUT_419F 16'h3BF1
`define CUBE_LUT_41A0 16'h3BF1
`define CUBE_LUT_41A1 16'h3BF1
`define CUBE_LUT_41A2 16'h3BF1
`define CUBE_LUT_41A3 16'h3BF1
`define CUBE_LUT_41A4 16'h3BF2
`define CUBE_LUT_41A5 16'h3BF2
`define CUBE_LUT_41A6 16'h3BF2
`define CUBE_LUT_41A7 16'h3BF2
`define CUBE_LUT_41A8 16'h3BF2
`define CUBE_LUT_41A9 16'h3BF2
`define CUBE_LUT_41AA 16'h3BF2
`define CUBE_LUT_41AB 16'h3BF2
`define CUBE_LUT_41AC 16'h3BF2
`define CUBE_LUT_41AD 16'h3BF2
`define CUBE_LUT_41AE 16'h3BF2
`define CUBE_LUT_41AF 16'h3BF2
`define CUBE_LUT_41B0 16'h3BF2
`define CUBE_LUT_41B1 16'h3BF2
`define CUBE_LUT_41B2 16'h3BF2
`define CUBE_LUT_41B3 16'h3BF2
`define CUBE_LUT_41B4 16'h3BF2
`define CUBE_LUT_41B5 16'h3BF2
`define CUBE_LUT_41B6 16'h3BF2
`define CUBE_LUT_41B7 16'h3BF3
`define CUBE_LUT_41B8 16'h3BF3
`define CUBE_LUT_41B9 16'h3BF3
`define CUBE_LUT_41BA 16'h3BF3
`define CUBE_LUT_41BB 16'h3BF3
`define CUBE_LUT_41BC 16'h3BF3
`define CUBE_LUT_41BD 16'h3BF3
`define CUBE_LUT_41BE 16'h3BF3
`define CUBE_LUT_41BF 16'h3BF3
`define CUBE_LUT_41C0 16'h3BF3
`define CUBE_LUT_41C1 16'h3BF3
`define CUBE_LUT_41C2 16'h3BF3
`define CUBE_LUT_41C3 16'h3BF3
`define CUBE_LUT_41C4 16'h3BF3
`define CUBE_LUT_41C5 16'h3BF3
`define CUBE_LUT_41C6 16'h3BF3
`define CUBE_LUT_41C7 16'h3BF3
`define CUBE_LUT_41C8 16'h3BF3
`define CUBE_LUT_41C9 16'h3BF3
`define CUBE_LUT_41CA 16'h3BF4
`define CUBE_LUT_41CB 16'h3BF4
`define CUBE_LUT_41CC 16'h3BF4
`define CUBE_LUT_41CD 16'h3BF4
`define CUBE_LUT_41CE 16'h3BF4
`define CUBE_LUT_41CF 16'h3BF4
`define CUBE_LUT_41D0 16'h3BF4
`define CUBE_LUT_41D1 16'h3BF4
`define CUBE_LUT_41D2 16'h3BF4
`define CUBE_LUT_41D3 16'h3BF4
`define CUBE_LUT_41D4 16'h3BF4
`define CUBE_LUT_41D5 16'h3BF4
`define CUBE_LUT_41D6 16'h3BF4
`define CUBE_LUT_41D7 16'h3BF4
`define CUBE_LUT_41D8 16'h3BF4
`define CUBE_LUT_41D9 16'h3BF4
`define CUBE_LUT_41DA 16'h3BF4
`define CUBE_LUT_41DB 16'h3BF4
`define CUBE_LUT_41DC 16'h3BF4
`define CUBE_LUT_41DD 16'h3BF4
`define CUBE_LUT_41DE 16'h3BF4
`define CUBE_LUT_41DF 16'h3BF4
`define CUBE_LUT_41E0 16'h3BF5
`define CUBE_LUT_41E1 16'h3BF5
`define CUBE_LUT_41E2 16'h3BF5
`define CUBE_LUT_41E3 16'h3BF5
`define CUBE_LUT_41E4 16'h3BF5
`define CUBE_LUT_41E5 16'h3BF5
`define CUBE_LUT_41E6 16'h3BF5
`define CUBE_LUT_41E7 16'h3BF5
`define CUBE_LUT_41E8 16'h3BF5
`define CUBE_LUT_41E9 16'h3BF5
`define CUBE_LUT_41EA 16'h3BF5
`define CUBE_LUT_41EB 16'h3BF5
`define CUBE_LUT_41EC 16'h3BF5
`define CUBE_LUT_41ED 16'h3BF5
`define CUBE_LUT_41EE 16'h3BF5
`define CUBE_LUT_41EF 16'h3BF5
`define CUBE_LUT_41F0 16'h3BF5
`define CUBE_LUT_41F1 16'h3BF5
`define CUBE_LUT_41F2 16'h3BF5
`define CUBE_LUT_41F3 16'h3BF5
`define CUBE_LUT_41F4 16'h3BF5
`define CUBE_LUT_41F5 16'h3BF5
`define CUBE_LUT_41F6 16'h3BF5
`define CUBE_LUT_41F7 16'h3BF6
`define CUBE_LUT_41F8 16'h3BF6
`define CUBE_LUT_41F9 16'h3BF6
`define CUBE_LUT_41FA 16'h3BF6
`define CUBE_LUT_41FB 16'h3BF6
`define CUBE_LUT_41FC 16'h3BF6
`define CUBE_LUT_41FD 16'h3BF6
`define CUBE_LUT_41FE 16'h3BF6
`define CUBE_LUT_41FF 16'h3BF6
`define CUBE_LUT_4200 16'h3BF6

`define CUBE_LUT_A895 16'hA894
`define CUBE_LUT_A896 16'hA895
`define CUBE_LUT_A897 16'hA896
`define CUBE_LUT_A898 16'hA897
`define CUBE_LUT_A899 16'hA898
`define CUBE_LUT_A89A 16'hA899
`define CUBE_LUT_A89B 16'hA89A
`define CUBE_LUT_A89C 16'hA89B
`define CUBE_LUT_A89D 16'hA89C
`define CUBE_LUT_A89E 16'hA89D
`define CUBE_LUT_A89F 16'hA89E
`define CUBE_LUT_A8A0 16'hA89F
`define CUBE_LUT_A8A1 16'hA8A0
`define CUBE_LUT_A8A2 16'hA8A1
`define CUBE_LUT_A8A3 16'hA8A2
`define CUBE_LUT_A8A4 16'hA8A3
`define CUBE_LUT_A8A5 16'hA8A4
`define CUBE_LUT_A8A6 16'hA8A5
`define CUBE_LUT_A8A7 16'hA8A6
`define CUBE_LUT_A8A8 16'hA8A7
`define CUBE_LUT_A8A9 16'hA8A8
`define CUBE_LUT_A8AA 16'hA8A9
`define CUBE_LUT_A8AB 16'hA8AA
`define CUBE_LUT_A8AC 16'hA8AB
`define CUBE_LUT_A8AD 16'hA8AC
`define CUBE_LUT_A8AE 16'hA8AD
`define CUBE_LUT_A8AF 16'hA8AE
`define CUBE_LUT_A8B0 16'hA8AF
`define CUBE_LUT_A8B1 16'hA8B0
`define CUBE_LUT_A8B2 16'hA8B1
`define CUBE_LUT_A8B3 16'hA8B2
`define CUBE_LUT_A8B4 16'hA8B3
`define CUBE_LUT_A8B5 16'hA8B4
`define CUBE_LUT_A8B6 16'hA8B5
`define CUBE_LUT_A8B7 16'hA8B6
`define CUBE_LUT_A8B8 16'hA8B7
`define CUBE_LUT_A8B9 16'hA8B8
`define CUBE_LUT_A8BA 16'hA8B9
`define CUBE_LUT_A8BB 16'hA8BA
`define CUBE_LUT_A8BC 16'hA8BB
`define CUBE_LUT_A8BD 16'hA8BC
`define CUBE_LUT_A8BE 16'hA8BD
`define CUBE_LUT_A8BF 16'hA8BE
`define CUBE_LUT_A8C0 16'hA8BF
`define CUBE_LUT_A8C1 16'hA8C0
`define CUBE_LUT_A8C2 16'hA8C1
`define CUBE_LUT_A8C3 16'hA8C2
`define CUBE_LUT_A8C4 16'hA8C3
`define CUBE_LUT_A8C5 16'hA8C4
`define CUBE_LUT_A8C6 16'hA8C5
`define CUBE_LUT_A8C7 16'hA8C6
`define CUBE_LUT_A8C8 16'hA8C7
`define CUBE_LUT_A8C9 16'hA8C8
`define CUBE_LUT_A8CA 16'hA8C9
`define CUBE_LUT_A8CB 16'hA8CA
`define CUBE_LUT_A8CC 16'hA8CB
`define CUBE_LUT_A8CD 16'hA8CC
`define CUBE_LUT_A8CE 16'hA8CD
`define CUBE_LUT_A8CF 16'hA8CE
`define CUBE_LUT_A8D0 16'hA8CF
`define CUBE_LUT_A8D1 16'hA8D0
`define CUBE_LUT_A8D2 16'hA8D1
`define CUBE_LUT_A8D3 16'hA8D2
`define CUBE_LUT_A8D4 16'hA8D3
`define CUBE_LUT_A8D5 16'hA8D4
`define CUBE_LUT_A8D6 16'hA8D5
`define CUBE_LUT_A8D7 16'hA8D6
`define CUBE_LUT_A8D8 16'hA8D7
`define CUBE_LUT_A8D9 16'hA8D8
`define CUBE_LUT_A8DA 16'hA8D9
`define CUBE_LUT_A8DB 16'hA8DA
`define CUBE_LUT_A8DC 16'hA8DB
`define CUBE_LUT_A8DD 16'hA8DC
`define CUBE_LUT_A8DE 16'hA8DD
`define CUBE_LUT_A8DF 16'hA8DE
`define CUBE_LUT_A8E0 16'hA8DF
`define CUBE_LUT_A8E1 16'hA8E0
`define CUBE_LUT_A8E2 16'hA8E1
`define CUBE_LUT_A8E3 16'hA8E2
`define CUBE_LUT_A8E4 16'hA8E3
`define CUBE_LUT_A8E5 16'hA8E4
`define CUBE_LUT_A8E6 16'hA8E5
`define CUBE_LUT_A8E7 16'hA8E6
`define CUBE_LUT_A8E8 16'hA8E7
`define CUBE_LUT_A8E9 16'hA8E8
`define CUBE_LUT_A8EA 16'hA8E9
`define CUBE_LUT_A8EB 16'hA8EA
`define CUBE_LUT_A8EC 16'hA8EB
`define CUBE_LUT_A8ED 16'hA8EC
`define CUBE_LUT_A8EE 16'hA8ED
`define CUBE_LUT_A8EF 16'hA8EE
`define CUBE_LUT_A8F0 16'hA8EF
`define CUBE_LUT_A8F1 16'hA8F0
`define CUBE_LUT_A8F2 16'hA8F1
`define CUBE_LUT_A8F3 16'hA8F2
`define CUBE_LUT_A8F4 16'hA8F3
`define CUBE_LUT_A8F5 16'hA8F4
`define CUBE_LUT_A8F6 16'hA8F5
`define CUBE_LUT_A8F7 16'hA8F6
`define CUBE_LUT_A8F8 16'hA8F7
`define CUBE_LUT_A8F9 16'hA8F8
`define CUBE_LUT_A8FA 16'hA8F9
`define CUBE_LUT_A8FB 16'hA8FA
`define CUBE_LUT_A8FC 16'hA8FB
`define CUBE_LUT_A8FD 16'hA8FC
`define CUBE_LUT_A8FE 16'hA8FD
`define CUBE_LUT_A8FF 16'hA8FE
`define CUBE_LUT_A900 16'hA8FF
`define CUBE_LUT_A901 16'hA900
`define CUBE_LUT_A902 16'hA901
`define CUBE_LUT_A903 16'hA902
`define CUBE_LUT_A904 16'hA903
`define CUBE_LUT_A905 16'hA904
`define CUBE_LUT_A906 16'hA905
`define CUBE_LUT_A907 16'hA906
`define CUBE_LUT_A908 16'hA907
`define CUBE_LUT_A909 16'hA908
`define CUBE_LUT_A90A 16'hA909
`define CUBE_LUT_A90B 16'hA90A
`define CUBE_LUT_A90C 16'hA90B
`define CUBE_LUT_A90D 16'hA90C
`define CUBE_LUT_A90E 16'hA90D
`define CUBE_LUT_A90F 16'hA90E
`define CUBE_LUT_A910 16'hA90F
`define CUBE_LUT_A911 16'hA910
`define CUBE_LUT_A912 16'hA911
`define CUBE_LUT_A913 16'hA912
`define CUBE_LUT_A914 16'hA913
`define CUBE_LUT_A915 16'hA914
`define CUBE_LUT_A916 16'hA915
`define CUBE_LUT_A917 16'hA916
`define CUBE_LUT_A918 16'hA917
`define CUBE_LUT_A919 16'hA918
`define CUBE_LUT_A91A 16'hA919
`define CUBE_LUT_A91B 16'hA91A
`define CUBE_LUT_A91C 16'hA91B
`define CUBE_LUT_A91D 16'hA91C
`define CUBE_LUT_A91E 16'hA91D
`define CUBE_LUT_A91F 16'hA91E
`define CUBE_LUT_A920 16'hA91F
`define CUBE_LUT_A921 16'hA920
`define CUBE_LUT_A922 16'hA921
`define CUBE_LUT_A923 16'hA922
`define CUBE_LUT_A924 16'hA923
`define CUBE_LUT_A925 16'hA924
`define CUBE_LUT_A926 16'hA925
`define CUBE_LUT_A927 16'hA926
`define CUBE_LUT_A928 16'hA927
`define CUBE_LUT_A929 16'hA928
`define CUBE_LUT_A92A 16'hA929
`define CUBE_LUT_A92B 16'hA92A
`define CUBE_LUT_A92C 16'hA92B
`define CUBE_LUT_A92D 16'hA92C
`define CUBE_LUT_A92E 16'hA92D
`define CUBE_LUT_A92F 16'hA92E
`define CUBE_LUT_A930 16'hA92F
`define CUBE_LUT_A931 16'hA930
`define CUBE_LUT_A932 16'hA931
`define CUBE_LUT_A933 16'hA932
`define CUBE_LUT_A934 16'hA933
`define CUBE_LUT_A935 16'hA934
`define CUBE_LUT_A936 16'hA935
`define CUBE_LUT_A937 16'hA936
`define CUBE_LUT_A938 16'hA937
`define CUBE_LUT_A939 16'hA938
`define CUBE_LUT_A93A 16'hA939
`define CUBE_LUT_A93B 16'hA93A
`define CUBE_LUT_A93C 16'hA93B
`define CUBE_LUT_A93D 16'hA93C
`define CUBE_LUT_A93E 16'hA93D
`define CUBE_LUT_A93F 16'hA93E
`define CUBE_LUT_A940 16'hA93F
`define CUBE_LUT_A941 16'hA940
`define CUBE_LUT_A942 16'hA941
`define CUBE_LUT_A943 16'hA942
`define CUBE_LUT_A944 16'hA943
`define CUBE_LUT_A945 16'hA944
`define CUBE_LUT_A946 16'hA945
`define CUBE_LUT_A947 16'hA946
`define CUBE_LUT_A948 16'hA947
`define CUBE_LUT_A949 16'hA948
`define CUBE_LUT_A94A 16'hA949
`define CUBE_LUT_A94B 16'hA94A
`define CUBE_LUT_A94C 16'hA94B
`define CUBE_LUT_A94D 16'hA94C
`define CUBE_LUT_A94E 16'hA94D
`define CUBE_LUT_A94F 16'hA94E
`define CUBE_LUT_A950 16'hA94F
`define CUBE_LUT_A951 16'hA950
`define CUBE_LUT_A952 16'hA951
`define CUBE_LUT_A953 16'hA952
`define CUBE_LUT_A954 16'hA953
`define CUBE_LUT_A955 16'hA954
`define CUBE_LUT_A956 16'hA955
`define CUBE_LUT_A957 16'hA956
`define CUBE_LUT_A958 16'hA957
`define CUBE_LUT_A959 16'hA958
`define CUBE_LUT_A95A 16'hA959
`define CUBE_LUT_A95B 16'hA95A
`define CUBE_LUT_A95C 16'hA95B
`define CUBE_LUT_A95D 16'hA95C
`define CUBE_LUT_A95E 16'hA95D
`define CUBE_LUT_A95F 16'hA95E
`define CUBE_LUT_A960 16'hA95F
`define CUBE_LUT_A961 16'hA960
`define CUBE_LUT_A962 16'hA961
`define CUBE_LUT_A963 16'hA962
`define CUBE_LUT_A964 16'hA963
`define CUBE_LUT_A965 16'hA964
`define CUBE_LUT_A966 16'hA965
`define CUBE_LUT_A967 16'hA966
`define CUBE_LUT_A968 16'hA967
`define CUBE_LUT_A969 16'hA968
`define CUBE_LUT_A96A 16'hA969
`define CUBE_LUT_A96B 16'hA96A
`define CUBE_LUT_A96C 16'hA96B
`define CUBE_LUT_A96D 16'hA96C
`define CUBE_LUT_A96E 16'hA96D
`define CUBE_LUT_A96F 16'hA96E
`define CUBE_LUT_A970 16'hA96F
`define CUBE_LUT_A971 16'hA970
`define CUBE_LUT_A972 16'hA971
`define CUBE_LUT_A973 16'hA972
`define CUBE_LUT_A974 16'hA973
`define CUBE_LUT_A975 16'hA974
`define CUBE_LUT_A976 16'hA975
`define CUBE_LUT_A977 16'hA976
`define CUBE_LUT_A978 16'hA977
`define CUBE_LUT_A979 16'hA978
`define CUBE_LUT_A97A 16'hA979
`define CUBE_LUT_A97B 16'hA97A
`define CUBE_LUT_A97C 16'hA97B
`define CUBE_LUT_A97D 16'hA97C
`define CUBE_LUT_A97E 16'hA97D
`define CUBE_LUT_A97F 16'hA97E
`define CUBE_LUT_A980 16'hA97F
`define CUBE_LUT_A981 16'hA980
`define CUBE_LUT_A982 16'hA981
`define CUBE_LUT_A983 16'hA982
`define CUBE_LUT_A984 16'hA983
`define CUBE_LUT_A985 16'hA984
`define CUBE_LUT_A986 16'hA985
`define CUBE_LUT_A987 16'hA986
`define CUBE_LUT_A988 16'hA987
`define CUBE_LUT_A989 16'hA988
`define CUBE_LUT_A98A 16'hA989
`define CUBE_LUT_A98B 16'hA98A
`define CUBE_LUT_A98C 16'hA98B
`define CUBE_LUT_A98D 16'hA98C
`define CUBE_LUT_A98E 16'hA98D
`define CUBE_LUT_A98F 16'hA98E
`define CUBE_LUT_A990 16'hA98F
`define CUBE_LUT_A991 16'hA990
`define CUBE_LUT_A992 16'hA991
`define CUBE_LUT_A993 16'hA992
`define CUBE_LUT_A994 16'hA993
`define CUBE_LUT_A995 16'hA994
`define CUBE_LUT_A996 16'hA995
`define CUBE_LUT_A997 16'hA996
`define CUBE_LUT_A998 16'hA997
`define CUBE_LUT_A999 16'hA998
`define CUBE_LUT_A99A 16'hA999
`define CUBE_LUT_A99B 16'hA99A
`define CUBE_LUT_A99C 16'hA99B
`define CUBE_LUT_A99D 16'hA99C
`define CUBE_LUT_A99E 16'hA99D
`define CUBE_LUT_A99F 16'hA99E
`define CUBE_LUT_A9A0 16'hA99F
`define CUBE_LUT_A9A1 16'hA9A0
`define CUBE_LUT_A9A2 16'hA9A1
`define CUBE_LUT_A9A3 16'hA9A2
`define CUBE_LUT_A9A4 16'hA9A3
`define CUBE_LUT_A9A5 16'hA9A4
`define CUBE_LUT_A9A6 16'hA9A5
`define CUBE_LUT_A9A7 16'hA9A6
`define CUBE_LUT_A9A8 16'hA9A7
`define CUBE_LUT_A9A9 16'hA9A8
`define CUBE_LUT_A9AA 16'hA9A9
`define CUBE_LUT_A9AB 16'hA9AA
`define CUBE_LUT_A9AC 16'hA9AB
`define CUBE_LUT_A9AD 16'hA9AC
`define CUBE_LUT_A9AE 16'hA9AD
`define CUBE_LUT_A9AF 16'hA9AE
`define CUBE_LUT_A9B0 16'hA9AF
`define CUBE_LUT_A9B1 16'hA9B0
`define CUBE_LUT_A9B2 16'hA9B1
`define CUBE_LUT_A9B3 16'hA9B2
`define CUBE_LUT_A9B4 16'hA9B3
`define CUBE_LUT_A9B5 16'hA9B4
`define CUBE_LUT_A9B6 16'hA9B5
`define CUBE_LUT_A9B7 16'hA9B6
`define CUBE_LUT_A9B8 16'hA9B7
`define CUBE_LUT_A9B9 16'hA9B8
`define CUBE_LUT_A9BA 16'hA9B9
`define CUBE_LUT_A9BB 16'hA9BA
`define CUBE_LUT_A9BC 16'hA9BB
`define CUBE_LUT_A9BD 16'hA9BC
`define CUBE_LUT_A9BE 16'hA9BD
`define CUBE_LUT_A9BF 16'hA9BE
`define CUBE_LUT_A9C0 16'hA9BF
`define CUBE_LUT_A9C1 16'hA9C0
`define CUBE_LUT_A9C2 16'hA9C1
`define CUBE_LUT_A9C3 16'hA9C2
`define CUBE_LUT_A9C4 16'hA9C3
`define CUBE_LUT_A9C5 16'hA9C4
`define CUBE_LUT_A9C6 16'hA9C5
`define CUBE_LUT_A9C7 16'hA9C6
`define CUBE_LUT_A9C8 16'hA9C7
`define CUBE_LUT_A9C9 16'hA9C8
`define CUBE_LUT_A9CA 16'hA9C9
`define CUBE_LUT_A9CB 16'hA9CA
`define CUBE_LUT_A9CC 16'hA9CB
`define CUBE_LUT_A9CD 16'hA9CC
`define CUBE_LUT_A9CE 16'hA9CD
`define CUBE_LUT_A9CF 16'hA9CE
`define CUBE_LUT_A9D0 16'hA9CF
`define CUBE_LUT_A9D1 16'hA9D0
`define CUBE_LUT_A9D2 16'hA9D1
`define CUBE_LUT_A9D3 16'hA9D2
`define CUBE_LUT_A9D4 16'hA9D3
`define CUBE_LUT_A9D5 16'hA9D4
`define CUBE_LUT_A9D6 16'hA9D5
`define CUBE_LUT_A9D7 16'hA9D6
`define CUBE_LUT_A9D8 16'hA9D7
`define CUBE_LUT_A9D9 16'hA9D8
`define CUBE_LUT_A9DA 16'hA9D9
`define CUBE_LUT_A9DB 16'hA9DA
`define CUBE_LUT_A9DC 16'hA9DB
`define CUBE_LUT_A9DD 16'hA9DC
`define CUBE_LUT_A9DE 16'hA9DD
`define CUBE_LUT_A9DF 16'hA9DE
`define CUBE_LUT_A9E0 16'hA9DF
`define CUBE_LUT_A9E1 16'hA9E0
`define CUBE_LUT_A9E2 16'hA9E1
`define CUBE_LUT_A9E3 16'hA9E2
`define CUBE_LUT_A9E4 16'hA9E3
`define CUBE_LUT_A9E5 16'hA9E4
`define CUBE_LUT_A9E6 16'hA9E5
`define CUBE_LUT_A9E7 16'hA9E6
`define CUBE_LUT_A9E8 16'hA9E7
`define CUBE_LUT_A9E9 16'hA9E8
`define CUBE_LUT_A9EA 16'hA9E9
`define CUBE_LUT_A9EB 16'hA9EA
`define CUBE_LUT_A9EC 16'hA9EB
`define CUBE_LUT_A9ED 16'hA9EC
`define CUBE_LUT_A9EE 16'hA9ED
`define CUBE_LUT_A9EF 16'hA9EE
`define CUBE_LUT_A9F0 16'hA9EF
`define CUBE_LUT_A9F1 16'hA9F0
`define CUBE_LUT_A9F2 16'hA9F1
`define CUBE_LUT_A9F3 16'hA9F2
`define CUBE_LUT_A9F4 16'hA9F3
`define CUBE_LUT_A9F5 16'hA9F4
`define CUBE_LUT_A9F6 16'hA9F5
`define CUBE_LUT_A9F7 16'hA9F6
`define CUBE_LUT_A9F8 16'hA9F7
`define CUBE_LUT_A9F9 16'hA9F8
`define CUBE_LUT_A9FA 16'hA9F9
`define CUBE_LUT_A9FB 16'hA9FA
`define CUBE_LUT_A9FC 16'hA9FB
`define CUBE_LUT_A9FD 16'hA9FC
`define CUBE_LUT_A9FE 16'hA9FD
`define CUBE_LUT_A9FF 16'hA9FE
`define CUBE_LUT_AA00 16'hA9FF
`define CUBE_LUT_AA01 16'hAA00
`define CUBE_LUT_AA02 16'hAA01
`define CUBE_LUT_AA03 16'hAA02
`define CUBE_LUT_AA04 16'hAA03
`define CUBE_LUT_AA05 16'hAA04
`define CUBE_LUT_AA06 16'hAA05
`define CUBE_LUT_AA07 16'hAA06
`define CUBE_LUT_AA08 16'hAA07
`define CUBE_LUT_AA09 16'hAA08
`define CUBE_LUT_AA0A 16'hAA09
`define CUBE_LUT_AA0B 16'hAA0A
`define CUBE_LUT_AA0C 16'hAA0B
`define CUBE_LUT_AA0D 16'hAA0C
`define CUBE_LUT_AA0E 16'hAA0D
`define CUBE_LUT_AA0F 16'hAA0E
`define CUBE_LUT_AA10 16'hAA0F
`define CUBE_LUT_AA11 16'hAA10
`define CUBE_LUT_AA12 16'hAA11
`define CUBE_LUT_AA13 16'hAA12
`define CUBE_LUT_AA14 16'hAA13
`define CUBE_LUT_AA15 16'hAA14
`define CUBE_LUT_AA16 16'hAA15
`define CUBE_LUT_AA17 16'hAA16
`define CUBE_LUT_AA18 16'hAA17
`define CUBE_LUT_AA19 16'hAA18
`define CUBE_LUT_AA1A 16'hAA19
`define CUBE_LUT_AA1B 16'hAA1A
`define CUBE_LUT_AA1C 16'hAA1B
`define CUBE_LUT_AA1D 16'hAA1C
`define CUBE_LUT_AA1E 16'hAA1D
`define CUBE_LUT_AA1F 16'hAA1E
`define CUBE_LUT_AA20 16'hAA1F
`define CUBE_LUT_AA21 16'hAA20
`define CUBE_LUT_AA22 16'hAA21
`define CUBE_LUT_AA23 16'hAA22
`define CUBE_LUT_AA24 16'hAA23
`define CUBE_LUT_AA25 16'hAA24
`define CUBE_LUT_AA26 16'hAA25
`define CUBE_LUT_AA27 16'hAA26
`define CUBE_LUT_AA28 16'hAA27
`define CUBE_LUT_AA29 16'hAA28
`define CUBE_LUT_AA2A 16'hAA29
`define CUBE_LUT_AA2B 16'hAA2A
`define CUBE_LUT_AA2C 16'hAA2B
`define CUBE_LUT_AA2D 16'hAA2C
`define CUBE_LUT_AA2E 16'hAA2D
`define CUBE_LUT_AA2F 16'hAA2E
`define CUBE_LUT_AA30 16'hAA2F
`define CUBE_LUT_AA31 16'hAA30
`define CUBE_LUT_AA32 16'hAA31
`define CUBE_LUT_AA33 16'hAA32
`define CUBE_LUT_AA34 16'hAA33
`define CUBE_LUT_AA35 16'hAA34
`define CUBE_LUT_AA36 16'hAA35
`define CUBE_LUT_AA37 16'hAA36
`define CUBE_LUT_AA38 16'hAA37
`define CUBE_LUT_AA39 16'hAA38
`define CUBE_LUT_AA3A 16'hAA39
`define CUBE_LUT_AA3B 16'hAA3A
`define CUBE_LUT_AA3C 16'hAA3B
`define CUBE_LUT_AA3D 16'hAA3C
`define CUBE_LUT_AA3E 16'hAA3D
`define CUBE_LUT_AA3F 16'hAA3E
`define CUBE_LUT_AA40 16'hAA3F
`define CUBE_LUT_AA41 16'hAA40
`define CUBE_LUT_AA42 16'hAA41
`define CUBE_LUT_AA43 16'hAA42
`define CUBE_LUT_AA44 16'hAA43
`define CUBE_LUT_AA45 16'hAA44
`define CUBE_LUT_AA46 16'hAA45
`define CUBE_LUT_AA47 16'hAA46
`define CUBE_LUT_AA48 16'hAA47
`define CUBE_LUT_AA49 16'hAA48
`define CUBE_LUT_AA4A 16'hAA49
`define CUBE_LUT_AA4B 16'hAA4A
`define CUBE_LUT_AA4C 16'hAA4B
`define CUBE_LUT_AA4D 16'hAA4C
`define CUBE_LUT_AA4E 16'hAA4D
`define CUBE_LUT_AA4F 16'hAA4E
`define CUBE_LUT_AA50 16'hAA4F
`define CUBE_LUT_AA51 16'hAA50
`define CUBE_LUT_AA52 16'hAA51
`define CUBE_LUT_AA53 16'hAA52
`define CUBE_LUT_AA54 16'hAA53
`define CUBE_LUT_AA55 16'hAA54
`define CUBE_LUT_AA56 16'hAA55
`define CUBE_LUT_AA57 16'hAA56
`define CUBE_LUT_AA58 16'hAA57
`define CUBE_LUT_AA59 16'hAA58
`define CUBE_LUT_AA5A 16'hAA59
`define CUBE_LUT_AA5B 16'hAA5A
`define CUBE_LUT_AA5C 16'hAA5B
`define CUBE_LUT_AA5D 16'hAA5C
`define CUBE_LUT_AA5E 16'hAA5D
`define CUBE_LUT_AA5F 16'hAA5E
`define CUBE_LUT_AA60 16'hAA5F
`define CUBE_LUT_AA61 16'hAA60
`define CUBE_LUT_AA62 16'hAA61
`define CUBE_LUT_AA63 16'hAA62
`define CUBE_LUT_AA64 16'hAA63
`define CUBE_LUT_AA65 16'hAA64
`define CUBE_LUT_AA66 16'hAA65
`define CUBE_LUT_AA67 16'hAA66
`define CUBE_LUT_AA68 16'hAA67
`define CUBE_LUT_AA69 16'hAA68
`define CUBE_LUT_AA6A 16'hAA69
`define CUBE_LUT_AA6B 16'hAA6A
`define CUBE_LUT_AA6C 16'hAA6B
`define CUBE_LUT_AA6D 16'hAA6C
`define CUBE_LUT_AA6E 16'hAA6D
`define CUBE_LUT_AA6F 16'hAA6E
`define CUBE_LUT_AA70 16'hAA6F
`define CUBE_LUT_AA71 16'hAA70
`define CUBE_LUT_AA72 16'hAA71
`define CUBE_LUT_AA73 16'hAA72
`define CUBE_LUT_AA74 16'hAA73
`define CUBE_LUT_AA75 16'hAA74
`define CUBE_LUT_AA76 16'hAA75
`define CUBE_LUT_AA77 16'hAA76
`define CUBE_LUT_AA78 16'hAA77
`define CUBE_LUT_AA79 16'hAA78
`define CUBE_LUT_AA7A 16'hAA79
`define CUBE_LUT_AA7B 16'hAA7A
`define CUBE_LUT_AA7C 16'hAA7B
`define CUBE_LUT_AA7D 16'hAA7C
`define CUBE_LUT_AA7E 16'hAA7D
`define CUBE_LUT_AA7F 16'hAA7E
`define CUBE_LUT_AA80 16'hAA7F
`define CUBE_LUT_AA81 16'hAA80
`define CUBE_LUT_AA82 16'hAA81
`define CUBE_LUT_AA83 16'hAA82
`define CUBE_LUT_AA84 16'hAA83
`define CUBE_LUT_AA85 16'hAA84
`define CUBE_LUT_AA86 16'hAA85
`define CUBE_LUT_AA87 16'hAA86
`define CUBE_LUT_AA88 16'hAA87
`define CUBE_LUT_AA89 16'hAA88
`define CUBE_LUT_AA8A 16'hAA89
`define CUBE_LUT_AA8B 16'hAA8A
`define CUBE_LUT_AA8C 16'hAA8B
`define CUBE_LUT_AA8D 16'hAA8C
`define CUBE_LUT_AA8E 16'hAA8D
`define CUBE_LUT_AA8F 16'hAA8E
`define CUBE_LUT_AA90 16'hAA8F
`define CUBE_LUT_AA91 16'hAA90
`define CUBE_LUT_AA92 16'hAA91
`define CUBE_LUT_AA93 16'hAA92
`define CUBE_LUT_AA94 16'hAA93
`define CUBE_LUT_AA95 16'hAA94
`define CUBE_LUT_AA96 16'hAA95
`define CUBE_LUT_AA97 16'hAA96
`define CUBE_LUT_AA98 16'hAA97
`define CUBE_LUT_AA99 16'hAA98
`define CUBE_LUT_AA9A 16'hAA99
`define CUBE_LUT_AA9B 16'hAA9A
`define CUBE_LUT_AA9C 16'hAA9A
`define CUBE_LUT_AA9D 16'hAA9B
`define CUBE_LUT_AA9E 16'hAA9C
`define CUBE_LUT_AA9F 16'hAA9D
`define CUBE_LUT_AAA0 16'hAA9E
`define CUBE_LUT_AAA1 16'hAA9F
`define CUBE_LUT_AAA2 16'hAAA0
`define CUBE_LUT_AAA3 16'hAAA1
`define CUBE_LUT_AAA4 16'hAAA2
`define CUBE_LUT_AAA5 16'hAAA3
`define CUBE_LUT_AAA6 16'hAAA4
`define CUBE_LUT_AAA7 16'hAAA5
`define CUBE_LUT_AAA8 16'hAAA6
`define CUBE_LUT_AAA9 16'hAAA7
`define CUBE_LUT_AAAA 16'hAAA8
`define CUBE_LUT_AAAB 16'hAAA9
`define CUBE_LUT_AAAC 16'hAAAA
`define CUBE_LUT_AAAD 16'hAAAB
`define CUBE_LUT_AAAE 16'hAAAC
`define CUBE_LUT_AAAF 16'hAAAD
`define CUBE_LUT_AAB0 16'hAAAE
`define CUBE_LUT_AAB1 16'hAAAF
`define CUBE_LUT_AAB2 16'hAAB0
`define CUBE_LUT_AAB3 16'hAAB1
`define CUBE_LUT_AAB4 16'hAAB2
`define CUBE_LUT_AAB5 16'hAAB3
`define CUBE_LUT_AAB6 16'hAAB4
`define CUBE_LUT_AAB7 16'hAAB5
`define CUBE_LUT_AAB8 16'hAAB6
`define CUBE_LUT_AAB9 16'hAAB7
`define CUBE_LUT_AABA 16'hAAB8
`define CUBE_LUT_AABB 16'hAAB9
`define CUBE_LUT_AABC 16'hAABA
`define CUBE_LUT_AABD 16'hAABB
`define CUBE_LUT_AABE 16'hAABC
`define CUBE_LUT_AABF 16'hAABD
`define CUBE_LUT_AAC0 16'hAABE
`define CUBE_LUT_AAC1 16'hAABF
`define CUBE_LUT_AAC2 16'hAAC0
`define CUBE_LUT_AAC3 16'hAAC1
`define CUBE_LUT_AAC4 16'hAAC2
`define CUBE_LUT_AAC5 16'hAAC3
`define CUBE_LUT_AAC6 16'hAAC4
`define CUBE_LUT_AAC7 16'hAAC5
`define CUBE_LUT_AAC8 16'hAAC6
`define CUBE_LUT_AAC9 16'hAAC7
`define CUBE_LUT_AACA 16'hAAC8
`define CUBE_LUT_AACB 16'hAAC9
`define CUBE_LUT_AACC 16'hAACA
`define CUBE_LUT_AACD 16'hAACB
`define CUBE_LUT_AACE 16'hAACC
`define CUBE_LUT_AACF 16'hAACD
`define CUBE_LUT_AAD0 16'hAACE
`define CUBE_LUT_AAD1 16'hAACF
`define CUBE_LUT_AAD2 16'hAAD0
`define CUBE_LUT_AAD3 16'hAAD1
`define CUBE_LUT_AAD4 16'hAAD2
`define CUBE_LUT_AAD5 16'hAAD3
`define CUBE_LUT_AAD6 16'hAAD4
`define CUBE_LUT_AAD7 16'hAAD5
`define CUBE_LUT_AAD8 16'hAAD6
`define CUBE_LUT_AAD9 16'hAAD7
`define CUBE_LUT_AADA 16'hAAD8
`define CUBE_LUT_AADB 16'hAAD9
`define CUBE_LUT_AADC 16'hAADA
`define CUBE_LUT_AADD 16'hAADB
`define CUBE_LUT_AADE 16'hAADC
`define CUBE_LUT_AADF 16'hAADD
`define CUBE_LUT_AAE0 16'hAADE
`define CUBE_LUT_AAE1 16'hAADF
`define CUBE_LUT_AAE2 16'hAAE0
`define CUBE_LUT_AAE3 16'hAAE1
`define CUBE_LUT_AAE4 16'hAAE2
`define CUBE_LUT_AAE5 16'hAAE3
`define CUBE_LUT_AAE6 16'hAAE4
`define CUBE_LUT_AAE7 16'hAAE5
`define CUBE_LUT_AAE8 16'hAAE6
`define CUBE_LUT_AAE9 16'hAAE7
`define CUBE_LUT_AAEA 16'hAAE8
`define CUBE_LUT_AAEB 16'hAAE9
`define CUBE_LUT_AAEC 16'hAAEA
`define CUBE_LUT_AAED 16'hAAEB
`define CUBE_LUT_AAEE 16'hAAEC
`define CUBE_LUT_AAEF 16'hAAED
`define CUBE_LUT_AAF0 16'hAAEE
`define CUBE_LUT_AAF1 16'hAAEF
`define CUBE_LUT_AAF2 16'hAAF0
`define CUBE_LUT_AAF3 16'hAAF1
`define CUBE_LUT_AAF4 16'hAAF2
`define CUBE_LUT_AAF5 16'hAAF3
`define CUBE_LUT_AAF6 16'hAAF4
`define CUBE_LUT_AAF7 16'hAAF5
`define CUBE_LUT_AAF8 16'hAAF6
`define CUBE_LUT_AAF9 16'hAAF7
`define CUBE_LUT_AAFA 16'hAAF8
`define CUBE_LUT_AAFB 16'hAAF9
`define CUBE_LUT_AAFC 16'hAAFA
`define CUBE_LUT_AAFD 16'hAAFB
`define CUBE_LUT_AAFE 16'hAAFC
`define CUBE_LUT_AAFF 16'hAAFD
`define CUBE_LUT_AB00 16'hAAFE
`define CUBE_LUT_AB01 16'hAAFF
`define CUBE_LUT_AB02 16'hAB00
`define CUBE_LUT_AB03 16'hAB01
`define CUBE_LUT_AB04 16'hAB02
`define CUBE_LUT_AB05 16'hAB03
`define CUBE_LUT_AB06 16'hAB04
`define CUBE_LUT_AB07 16'hAB05
`define CUBE_LUT_AB08 16'hAB06
`define CUBE_LUT_AB09 16'hAB07
`define CUBE_LUT_AB0A 16'hAB08
`define CUBE_LUT_AB0B 16'hAB09
`define CUBE_LUT_AB0C 16'hAB0A
`define CUBE_LUT_AB0D 16'hAB0B
`define CUBE_LUT_AB0E 16'hAB0C
`define CUBE_LUT_AB0F 16'hAB0D
`define CUBE_LUT_AB10 16'hAB0E
`define CUBE_LUT_AB11 16'hAB0F
`define CUBE_LUT_AB12 16'hAB10
`define CUBE_LUT_AB13 16'hAB11
`define CUBE_LUT_AB14 16'hAB12
`define CUBE_LUT_AB15 16'hAB13
`define CUBE_LUT_AB16 16'hAB14
`define CUBE_LUT_AB17 16'hAB15
`define CUBE_LUT_AB18 16'hAB16
`define CUBE_LUT_AB19 16'hAB17
`define CUBE_LUT_AB1A 16'hAB18
`define CUBE_LUT_AB1B 16'hAB19
`define CUBE_LUT_AB1C 16'hAB1A
`define CUBE_LUT_AB1D 16'hAB1B
`define CUBE_LUT_AB1E 16'hAB1C
`define CUBE_LUT_AB1F 16'hAB1D
`define CUBE_LUT_AB20 16'hAB1E
`define CUBE_LUT_AB21 16'hAB1F
`define CUBE_LUT_AB22 16'hAB20
`define CUBE_LUT_AB23 16'hAB21
`define CUBE_LUT_AB24 16'hAB22
`define CUBE_LUT_AB25 16'hAB23
`define CUBE_LUT_AB26 16'hAB24
`define CUBE_LUT_AB27 16'hAB25
`define CUBE_LUT_AB28 16'hAB26
`define CUBE_LUT_AB29 16'hAB27
`define CUBE_LUT_AB2A 16'hAB28
`define CUBE_LUT_AB2B 16'hAB29
`define CUBE_LUT_AB2C 16'hAB2A
`define CUBE_LUT_AB2D 16'hAB2B
`define CUBE_LUT_AB2E 16'hAB2C
`define CUBE_LUT_AB2F 16'hAB2D
`define CUBE_LUT_AB30 16'hAB2E
`define CUBE_LUT_AB31 16'hAB2F
`define CUBE_LUT_AB32 16'hAB30
`define CUBE_LUT_AB33 16'hAB31
`define CUBE_LUT_AB34 16'hAB32
`define CUBE_LUT_AB35 16'hAB33
`define CUBE_LUT_AB36 16'hAB34
`define CUBE_LUT_AB37 16'hAB35
`define CUBE_LUT_AB38 16'hAB36
`define CUBE_LUT_AB39 16'hAB37
`define CUBE_LUT_AB3A 16'hAB38
`define CUBE_LUT_AB3B 16'hAB39
`define CUBE_LUT_AB3C 16'hAB3A
`define CUBE_LUT_AB3D 16'hAB3B
`define CUBE_LUT_AB3E 16'hAB3C
`define CUBE_LUT_AB3F 16'hAB3D
`define CUBE_LUT_AB40 16'hAB3E
`define CUBE_LUT_AB41 16'hAB3F
`define CUBE_LUT_AB42 16'hAB40
`define CUBE_LUT_AB43 16'hAB41
`define CUBE_LUT_AB44 16'hAB42
`define CUBE_LUT_AB45 16'hAB43
`define CUBE_LUT_AB46 16'hAB44
`define CUBE_LUT_AB47 16'hAB45
`define CUBE_LUT_AB48 16'hAB46
`define CUBE_LUT_AB49 16'hAB47
`define CUBE_LUT_AB4A 16'hAB48
`define CUBE_LUT_AB4B 16'hAB49
`define CUBE_LUT_AB4C 16'hAB4A
`define CUBE_LUT_AB4D 16'hAB4B
`define CUBE_LUT_AB4E 16'hAB4C
`define CUBE_LUT_AB4F 16'hAB4D
`define CUBE_LUT_AB50 16'hAB4E
`define CUBE_LUT_AB51 16'hAB4F
`define CUBE_LUT_AB52 16'hAB50
`define CUBE_LUT_AB53 16'hAB51
`define CUBE_LUT_AB54 16'hAB52
`define CUBE_LUT_AB55 16'hAB53
`define CUBE_LUT_AB56 16'hAB54
`define CUBE_LUT_AB57 16'hAB55
`define CUBE_LUT_AB58 16'hAB56
`define CUBE_LUT_AB59 16'hAB57
`define CUBE_LUT_AB5A 16'hAB58
`define CUBE_LUT_AB5B 16'hAB59
`define CUBE_LUT_AB5C 16'hAB5A
`define CUBE_LUT_AB5D 16'hAB5B
`define CUBE_LUT_AB5E 16'hAB5C
`define CUBE_LUT_AB5F 16'hAB5D
`define CUBE_LUT_AB60 16'hAB5E
`define CUBE_LUT_AB61 16'hAB5F
`define CUBE_LUT_AB62 16'hAB60
`define CUBE_LUT_AB63 16'hAB61
`define CUBE_LUT_AB64 16'hAB62
`define CUBE_LUT_AB65 16'hAB63
`define CUBE_LUT_AB66 16'hAB64
`define CUBE_LUT_AB67 16'hAB65
`define CUBE_LUT_AB68 16'hAB66
`define CUBE_LUT_AB69 16'hAB67
`define CUBE_LUT_AB6A 16'hAB68
`define CUBE_LUT_AB6B 16'hAB69
`define CUBE_LUT_AB6C 16'hAB6A
`define CUBE_LUT_AB6D 16'hAB6B
`define CUBE_LUT_AB6E 16'hAB6C
`define CUBE_LUT_AB6F 16'hAB6D
`define CUBE_LUT_AB70 16'hAB6E
`define CUBE_LUT_AB71 16'hAB6F
`define CUBE_LUT_AB72 16'hAB70
`define CUBE_LUT_AB73 16'hAB71
`define CUBE_LUT_AB74 16'hAB72
`define CUBE_LUT_AB75 16'hAB73
`define CUBE_LUT_AB76 16'hAB74
`define CUBE_LUT_AB77 16'hAB75
`define CUBE_LUT_AB78 16'hAB76
`define CUBE_LUT_AB79 16'hAB77
`define CUBE_LUT_AB7A 16'hAB78
`define CUBE_LUT_AB7B 16'hAB79
`define CUBE_LUT_AB7C 16'hAB7A
`define CUBE_LUT_AB7D 16'hAB7B
`define CUBE_LUT_AB7E 16'hAB7C
`define CUBE_LUT_AB7F 16'hAB7D
`define CUBE_LUT_AB80 16'hAB7E
`define CUBE_LUT_AB81 16'hAB7F
`define CUBE_LUT_AB82 16'hAB80
`define CUBE_LUT_AB83 16'hAB81
`define CUBE_LUT_AB84 16'hAB82
`define CUBE_LUT_AB85 16'hAB83
`define CUBE_LUT_AB86 16'hAB84
`define CUBE_LUT_AB87 16'hAB85
`define CUBE_LUT_AB88 16'hAB86
`define CUBE_LUT_AB89 16'hAB87
`define CUBE_LUT_AB8A 16'hAB88
`define CUBE_LUT_AB8B 16'hAB89
`define CUBE_LUT_AB8C 16'hAB8A
`define CUBE_LUT_AB8D 16'hAB8B
`define CUBE_LUT_AB8E 16'hAB8C
`define CUBE_LUT_AB8F 16'hAB8D
`define CUBE_LUT_AB90 16'hAB8E
`define CUBE_LUT_AB91 16'hAB8F
`define CUBE_LUT_AB92 16'hAB90
`define CUBE_LUT_AB93 16'hAB91
`define CUBE_LUT_AB94 16'hAB92
`define CUBE_LUT_AB95 16'hAB93
`define CUBE_LUT_AB96 16'hAB94
`define CUBE_LUT_AB97 16'hAB95
`define CUBE_LUT_AB98 16'hAB96
`define CUBE_LUT_AB99 16'hAB97
`define CUBE_LUT_AB9A 16'hAB98
`define CUBE_LUT_AB9B 16'hAB99
`define CUBE_LUT_AB9C 16'hAB9A
`define CUBE_LUT_AB9D 16'hAB9B
`define CUBE_LUT_AB9E 16'hAB9C
`define CUBE_LUT_AB9F 16'hAB9D
`define CUBE_LUT_ABA0 16'hAB9E
`define CUBE_LUT_ABA1 16'hAB9F
`define CUBE_LUT_ABA2 16'hABA0
`define CUBE_LUT_ABA3 16'hABA1
`define CUBE_LUT_ABA4 16'hABA2
`define CUBE_LUT_ABA5 16'hABA3
`define CUBE_LUT_ABA6 16'hABA4
`define CUBE_LUT_ABA7 16'hABA5
`define CUBE_LUT_ABA8 16'hABA6
`define CUBE_LUT_ABA9 16'hABA7
`define CUBE_LUT_ABAA 16'hABA8
`define CUBE_LUT_ABAB 16'hABA9
`define CUBE_LUT_ABAC 16'hABAA
`define CUBE_LUT_ABAD 16'hABAB
`define CUBE_LUT_ABAE 16'hABAC
`define CUBE_LUT_ABAF 16'hABAD
`define CUBE_LUT_ABB0 16'hABAE
`define CUBE_LUT_ABB1 16'hABAF
`define CUBE_LUT_ABB2 16'hABB0
`define CUBE_LUT_ABB3 16'hABB1
`define CUBE_LUT_ABB4 16'hABB2
`define CUBE_LUT_ABB5 16'hABB3
`define CUBE_LUT_ABB6 16'hABB4
`define CUBE_LUT_ABB7 16'hABB5
`define CUBE_LUT_ABB8 16'hABB6
`define CUBE_LUT_ABB9 16'hABB7
`define CUBE_LUT_ABBA 16'hABB8
`define CUBE_LUT_ABBB 16'hABB9
`define CUBE_LUT_ABBC 16'hABBA
`define CUBE_LUT_ABBD 16'hABBB
`define CUBE_LUT_ABBE 16'hABBC
`define CUBE_LUT_ABBF 16'hABBD
`define CUBE_LUT_ABC0 16'hABBE
`define CUBE_LUT_ABC1 16'hABBF
`define CUBE_LUT_ABC2 16'hABC0
`define CUBE_LUT_ABC3 16'hABC1
`define CUBE_LUT_ABC4 16'hABC2
`define CUBE_LUT_ABC5 16'hABC3
`define CUBE_LUT_ABC6 16'hABC4
`define CUBE_LUT_ABC7 16'hABC5
`define CUBE_LUT_ABC8 16'hABC6
`define CUBE_LUT_ABC9 16'hABC7
`define CUBE_LUT_ABCA 16'hABC8
`define CUBE_LUT_ABCB 16'hABC9
`define CUBE_LUT_ABCC 16'hABCA
`define CUBE_LUT_ABCD 16'hABCB
`define CUBE_LUT_ABCE 16'hABCC
`define CUBE_LUT_ABCF 16'hABCD
`define CUBE_LUT_ABD0 16'hABCE
`define CUBE_LUT_ABD1 16'hABCF
`define CUBE_LUT_ABD2 16'hABD0
`define CUBE_LUT_ABD3 16'hABD1
`define CUBE_LUT_ABD4 16'hABD2
`define CUBE_LUT_ABD5 16'hABD3
`define CUBE_LUT_ABD6 16'hABD3
`define CUBE_LUT_ABD7 16'hABD4
`define CUBE_LUT_ABD8 16'hABD5
`define CUBE_LUT_ABD9 16'hABD6
`define CUBE_LUT_ABDA 16'hABD7
`define CUBE_LUT_ABDB 16'hABD8
`define CUBE_LUT_ABDC 16'hABD9
`define CUBE_LUT_ABDD 16'hABDA
`define CUBE_LUT_ABDE 16'hABDB
`define CUBE_LUT_ABDF 16'hABDC
`define CUBE_LUT_ABE0 16'hABDD
`define CUBE_LUT_ABE1 16'hABDE
`define CUBE_LUT_ABE2 16'hABDF
`define CUBE_LUT_ABE3 16'hABE0
`define CUBE_LUT_ABE4 16'hABE1
`define CUBE_LUT_ABE5 16'hABE2
`define CUBE_LUT_ABE6 16'hABE3
`define CUBE_LUT_ABE7 16'hABE4
`define CUBE_LUT_ABE8 16'hABE5
`define CUBE_LUT_ABE9 16'hABE6
`define CUBE_LUT_ABEA 16'hABE7
`define CUBE_LUT_ABEB 16'hABE8
`define CUBE_LUT_ABEC 16'hABE9
`define CUBE_LUT_ABED 16'hABEA
`define CUBE_LUT_ABEE 16'hABEB
`define CUBE_LUT_ABEF 16'hABEC
`define CUBE_LUT_ABF0 16'hABED
`define CUBE_LUT_ABF1 16'hABEE
`define CUBE_LUT_ABF2 16'hABEF
`define CUBE_LUT_ABF3 16'hABF0
`define CUBE_LUT_ABF4 16'hABF1
`define CUBE_LUT_ABF5 16'hABF2
`define CUBE_LUT_ABF6 16'hABF3
`define CUBE_LUT_ABF7 16'hABF4
`define CUBE_LUT_ABF8 16'hABF5
`define CUBE_LUT_ABF9 16'hABF6
`define CUBE_LUT_ABFA 16'hABF7
`define CUBE_LUT_ABFB 16'hABF8
`define CUBE_LUT_ABFC 16'hABF9
`define CUBE_LUT_ABFD 16'hABFA
`define CUBE_LUT_ABFE 16'hABFB
`define CUBE_LUT_ABFF 16'hABFC
`define CUBE_LUT_AC00 16'hABFD
`define CUBE_LUT_AC01 16'hABFF
`define CUBE_LUT_AC02 16'hAC01
`define CUBE_LUT_AC03 16'hAC02
`define CUBE_LUT_AC04 16'hAC03
`define CUBE_LUT_AC05 16'hAC04
`define CUBE_LUT_AC06 16'hAC05
`define CUBE_LUT_AC07 16'hAC06
`define CUBE_LUT_AC08 16'hAC07
`define CUBE_LUT_AC09 16'hAC08
`define CUBE_LUT_AC0A 16'hAC09
`define CUBE_LUT_AC0B 16'hAC0A
`define CUBE_LUT_AC0C 16'hAC0B
`define CUBE_LUT_AC0D 16'hAC0C
`define CUBE_LUT_AC0E 16'hAC0D
`define CUBE_LUT_AC0F 16'hAC0E
`define CUBE_LUT_AC10 16'hAC0F
`define CUBE_LUT_AC11 16'hAC10
`define CUBE_LUT_AC12 16'hAC11
`define CUBE_LUT_AC13 16'hAC12
`define CUBE_LUT_AC14 16'hAC13
`define CUBE_LUT_AC15 16'hAC14
`define CUBE_LUT_AC16 16'hAC15
`define CUBE_LUT_AC17 16'hAC16
`define CUBE_LUT_AC18 16'hAC17
`define CUBE_LUT_AC19 16'hAC18
`define CUBE_LUT_AC1A 16'hAC19
`define CUBE_LUT_AC1B 16'hAC1A
`define CUBE_LUT_AC1C 16'hAC1B
`define CUBE_LUT_AC1D 16'hAC1C
`define CUBE_LUT_AC1E 16'hAC1D
`define CUBE_LUT_AC1F 16'hAC1E
`define CUBE_LUT_AC20 16'hAC1F
`define CUBE_LUT_AC21 16'hAC20
`define CUBE_LUT_AC22 16'hAC21
`define CUBE_LUT_AC23 16'hAC22
`define CUBE_LUT_AC24 16'hAC23
`define CUBE_LUT_AC25 16'hAC24
`define CUBE_LUT_AC26 16'hAC25
`define CUBE_LUT_AC27 16'hAC26
`define CUBE_LUT_AC28 16'hAC27
`define CUBE_LUT_AC29 16'hAC28
`define CUBE_LUT_AC2A 16'hAC28
`define CUBE_LUT_AC2B 16'hAC29
`define CUBE_LUT_AC2C 16'hAC2A
`define CUBE_LUT_AC2D 16'hAC2B
`define CUBE_LUT_AC2E 16'hAC2C
`define CUBE_LUT_AC2F 16'hAC2D
`define CUBE_LUT_AC30 16'hAC2E
`define CUBE_LUT_AC31 16'hAC2F
`define CUBE_LUT_AC32 16'hAC30
`define CUBE_LUT_AC33 16'hAC31
`define CUBE_LUT_AC34 16'hAC32
`define CUBE_LUT_AC35 16'hAC33
`define CUBE_LUT_AC36 16'hAC34
`define CUBE_LUT_AC37 16'hAC35
`define CUBE_LUT_AC38 16'hAC36
`define CUBE_LUT_AC39 16'hAC37
`define CUBE_LUT_AC3A 16'hAC38
`define CUBE_LUT_AC3B 16'hAC39
`define CUBE_LUT_AC3C 16'hAC3A
`define CUBE_LUT_AC3D 16'hAC3B
`define CUBE_LUT_AC3E 16'hAC3C
`define CUBE_LUT_AC3F 16'hAC3D
`define CUBE_LUT_AC40 16'hAC3E
`define CUBE_LUT_AC41 16'hAC3F
`define CUBE_LUT_AC42 16'hAC40
`define CUBE_LUT_AC43 16'hAC41
`define CUBE_LUT_AC44 16'hAC42
`define CUBE_LUT_AC45 16'hAC43
`define CUBE_LUT_AC46 16'hAC44
`define CUBE_LUT_AC47 16'hAC45
`define CUBE_LUT_AC48 16'hAC46
`define CUBE_LUT_AC49 16'hAC47
`define CUBE_LUT_AC4A 16'hAC48
`define CUBE_LUT_AC4B 16'hAC49
`define CUBE_LUT_AC4C 16'hAC4A
`define CUBE_LUT_AC4D 16'hAC4B
`define CUBE_LUT_AC4E 16'hAC4C
`define CUBE_LUT_AC4F 16'hAC4D
`define CUBE_LUT_AC50 16'hAC4E
`define CUBE_LUT_AC51 16'hAC4F
`define CUBE_LUT_AC52 16'hAC50
`define CUBE_LUT_AC53 16'hAC51
`define CUBE_LUT_AC54 16'hAC52
`define CUBE_LUT_AC55 16'hAC53
`define CUBE_LUT_AC56 16'hAC54
`define CUBE_LUT_AC57 16'hAC55
`define CUBE_LUT_AC58 16'hAC56
`define CUBE_LUT_AC59 16'hAC57
`define CUBE_LUT_AC5A 16'hAC58
`define CUBE_LUT_AC5B 16'hAC59
`define CUBE_LUT_AC5C 16'hAC5A
`define CUBE_LUT_AC5D 16'hAC5B
`define CUBE_LUT_AC5E 16'hAC5C
`define CUBE_LUT_AC5F 16'hAC5D
`define CUBE_LUT_AC60 16'hAC5E
`define CUBE_LUT_AC61 16'hAC5F
`define CUBE_LUT_AC62 16'hAC60
`define CUBE_LUT_AC63 16'hAC61
`define CUBE_LUT_AC64 16'hAC62
`define CUBE_LUT_AC65 16'hAC63
`define CUBE_LUT_AC66 16'hAC64
`define CUBE_LUT_AC67 16'hAC65
`define CUBE_LUT_AC68 16'hAC66
`define CUBE_LUT_AC69 16'hAC67
`define CUBE_LUT_AC6A 16'hAC68
`define CUBE_LUT_AC6B 16'hAC69
`define CUBE_LUT_AC6C 16'hAC6A
`define CUBE_LUT_AC6D 16'hAC6B
`define CUBE_LUT_AC6E 16'hAC6C
`define CUBE_LUT_AC6F 16'hAC6D
`define CUBE_LUT_AC70 16'hAC6E
`define CUBE_LUT_AC71 16'hAC6F
`define CUBE_LUT_AC72 16'hAC70
`define CUBE_LUT_AC73 16'hAC71
`define CUBE_LUT_AC74 16'hAC72
`define CUBE_LUT_AC75 16'hAC73
`define CUBE_LUT_AC76 16'hAC74
`define CUBE_LUT_AC77 16'hAC75
`define CUBE_LUT_AC78 16'hAC76
`define CUBE_LUT_AC79 16'hAC77
`define CUBE_LUT_AC7A 16'hAC78
`define CUBE_LUT_AC7B 16'hAC79
`define CUBE_LUT_AC7C 16'hAC7A
`define CUBE_LUT_AC7D 16'hAC7B
`define CUBE_LUT_AC7E 16'hAC7C
`define CUBE_LUT_AC7F 16'hAC7D
`define CUBE_LUT_AC80 16'hAC7E
`define CUBE_LUT_AC81 16'hAC7F
`define CUBE_LUT_AC82 16'hAC80
`define CUBE_LUT_AC83 16'hAC81
`define CUBE_LUT_AC84 16'hAC82
`define CUBE_LUT_AC85 16'hAC83
`define CUBE_LUT_AC86 16'hAC84
`define CUBE_LUT_AC87 16'hAC85
`define CUBE_LUT_AC88 16'hAC86
`define CUBE_LUT_AC89 16'hAC87
`define CUBE_LUT_AC8A 16'hAC88
`define CUBE_LUT_AC8B 16'hAC89
`define CUBE_LUT_AC8C 16'hAC8A
`define CUBE_LUT_AC8D 16'hAC8B
`define CUBE_LUT_AC8E 16'hAC8C
`define CUBE_LUT_AC8F 16'hAC8D
`define CUBE_LUT_AC90 16'hAC8E
`define CUBE_LUT_AC91 16'hAC8F
`define CUBE_LUT_AC92 16'hAC90
`define CUBE_LUT_AC93 16'hAC91
`define CUBE_LUT_AC94 16'hAC92
`define CUBE_LUT_AC95 16'hAC93
`define CUBE_LUT_AC96 16'hAC94
`define CUBE_LUT_AC97 16'hAC95
`define CUBE_LUT_AC98 16'hAC96
`define CUBE_LUT_AC99 16'hAC97
`define CUBE_LUT_AC9A 16'hAC98
`define CUBE_LUT_AC9B 16'hAC99
`define CUBE_LUT_AC9C 16'hAC9A
`define CUBE_LUT_AC9D 16'hAC9B
`define CUBE_LUT_AC9E 16'hAC9C
`define CUBE_LUT_AC9F 16'hAC9D
`define CUBE_LUT_ACA0 16'hAC9E
`define CUBE_LUT_ACA1 16'hAC9F
`define CUBE_LUT_ACA2 16'hACA0
`define CUBE_LUT_ACA3 16'hACA1
`define CUBE_LUT_ACA4 16'hACA2
`define CUBE_LUT_ACA5 16'hACA3
`define CUBE_LUT_ACA6 16'hACA4
`define CUBE_LUT_ACA7 16'hACA5
`define CUBE_LUT_ACA8 16'hACA6
`define CUBE_LUT_ACA9 16'hACA7
`define CUBE_LUT_ACAA 16'hACA8
`define CUBE_LUT_ACAB 16'hACA9
`define CUBE_LUT_ACAC 16'hACAA
`define CUBE_LUT_ACAD 16'hACAB
`define CUBE_LUT_ACAE 16'hACAC
`define CUBE_LUT_ACAF 16'hACAD
`define CUBE_LUT_ACB0 16'hACAE
`define CUBE_LUT_ACB1 16'hACAF
`define CUBE_LUT_ACB2 16'hACB0
`define CUBE_LUT_ACB3 16'hACB1
`define CUBE_LUT_ACB4 16'hACB2
`define CUBE_LUT_ACB5 16'hACB3
`define CUBE_LUT_ACB6 16'hACB4
`define CUBE_LUT_ACB7 16'hACB5
`define CUBE_LUT_ACB8 16'hACB6
`define CUBE_LUT_ACB9 16'hACB7
`define CUBE_LUT_ACBA 16'hACB8
`define CUBE_LUT_ACBB 16'hACB9
`define CUBE_LUT_ACBC 16'hACBA
`define CUBE_LUT_ACBD 16'hACBB
`define CUBE_LUT_ACBE 16'hACBC
`define CUBE_LUT_ACBF 16'hACBD
`define CUBE_LUT_ACC0 16'hACBE
`define CUBE_LUT_ACC1 16'hACBF
`define CUBE_LUT_ACC2 16'hACC0
`define CUBE_LUT_ACC3 16'hACC1
`define CUBE_LUT_ACC4 16'hACC2
`define CUBE_LUT_ACC5 16'hACC3
`define CUBE_LUT_ACC6 16'hACC4
`define CUBE_LUT_ACC7 16'hACC5
`define CUBE_LUT_ACC8 16'hACC6
`define CUBE_LUT_ACC9 16'hACC7
`define CUBE_LUT_ACCA 16'hACC8
`define CUBE_LUT_ACCB 16'hACC9
`define CUBE_LUT_ACCC 16'hACCA
`define CUBE_LUT_ACCD 16'hACCB
`define CUBE_LUT_ACCE 16'hACCC
`define CUBE_LUT_ACCF 16'hACCD
`define CUBE_LUT_ACD0 16'hACCE
`define CUBE_LUT_ACD1 16'hACCF
`define CUBE_LUT_ACD2 16'hACD0
`define CUBE_LUT_ACD3 16'hACD1
`define CUBE_LUT_ACD4 16'hACD2
`define CUBE_LUT_ACD5 16'hACD3
`define CUBE_LUT_ACD6 16'hACD4
`define CUBE_LUT_ACD7 16'hACD5
`define CUBE_LUT_ACD8 16'hACD6
`define CUBE_LUT_ACD9 16'hACD7
`define CUBE_LUT_ACDA 16'hACD8
`define CUBE_LUT_ACDB 16'hACD9
`define CUBE_LUT_ACDC 16'hACDA
`define CUBE_LUT_ACDD 16'hACDB
`define CUBE_LUT_ACDE 16'hACDC
`define CUBE_LUT_ACDF 16'hACDD
`define CUBE_LUT_ACE0 16'hACDE
`define CUBE_LUT_ACE1 16'hACDF
`define CUBE_LUT_ACE2 16'hACE0
`define CUBE_LUT_ACE3 16'hACE1
`define CUBE_LUT_ACE4 16'hACE2
`define CUBE_LUT_ACE5 16'hACE3
`define CUBE_LUT_ACE6 16'hACE4
`define CUBE_LUT_ACE7 16'hACE5
`define CUBE_LUT_ACE8 16'hACE6
`define CUBE_LUT_ACE9 16'hACE7
`define CUBE_LUT_ACEA 16'hACE8
`define CUBE_LUT_ACEB 16'hACE9
`define CUBE_LUT_ACEC 16'hACEA
`define CUBE_LUT_ACED 16'hACEB
`define CUBE_LUT_ACEE 16'hACEC
`define CUBE_LUT_ACEF 16'hACED
`define CUBE_LUT_ACF0 16'hACED
`define CUBE_LUT_ACF1 16'hACEE
`define CUBE_LUT_ACF2 16'hACEF
`define CUBE_LUT_ACF3 16'hACF0
`define CUBE_LUT_ACF4 16'hACF1
`define CUBE_LUT_ACF5 16'hACF2
`define CUBE_LUT_ACF6 16'hACF3
`define CUBE_LUT_ACF7 16'hACF4
`define CUBE_LUT_ACF8 16'hACF5
`define CUBE_LUT_ACF9 16'hACF6
`define CUBE_LUT_ACFA 16'hACF7
`define CUBE_LUT_ACFB 16'hACF8
`define CUBE_LUT_ACFC 16'hACF9
`define CUBE_LUT_ACFD 16'hACFA
`define CUBE_LUT_ACFE 16'hACFB
`define CUBE_LUT_ACFF 16'hACFC
`define CUBE_LUT_AD00 16'hACFD
`define CUBE_LUT_AD01 16'hACFE
`define CUBE_LUT_AD02 16'hACFF
`define CUBE_LUT_AD03 16'hAD00
`define CUBE_LUT_AD04 16'hAD01
`define CUBE_LUT_AD05 16'hAD02
`define CUBE_LUT_AD06 16'hAD03
`define CUBE_LUT_AD07 16'hAD04
`define CUBE_LUT_AD08 16'hAD05
`define CUBE_LUT_AD09 16'hAD06
`define CUBE_LUT_AD0A 16'hAD07
`define CUBE_LUT_AD0B 16'hAD08
`define CUBE_LUT_AD0C 16'hAD09
`define CUBE_LUT_AD0D 16'hAD0A
`define CUBE_LUT_AD0E 16'hAD0B
`define CUBE_LUT_AD0F 16'hAD0C
`define CUBE_LUT_AD10 16'hAD0D
`define CUBE_LUT_AD11 16'hAD0E
`define CUBE_LUT_AD12 16'hAD0F
`define CUBE_LUT_AD13 16'hAD10
`define CUBE_LUT_AD14 16'hAD11
`define CUBE_LUT_AD15 16'hAD12
`define CUBE_LUT_AD16 16'hAD13
`define CUBE_LUT_AD17 16'hAD14
`define CUBE_LUT_AD18 16'hAD15
`define CUBE_LUT_AD19 16'hAD16
`define CUBE_LUT_AD1A 16'hAD17
`define CUBE_LUT_AD1B 16'hAD18
`define CUBE_LUT_AD1C 16'hAD19
`define CUBE_LUT_AD1D 16'hAD1A
`define CUBE_LUT_AD1E 16'hAD1B
`define CUBE_LUT_AD1F 16'hAD1C
`define CUBE_LUT_AD20 16'hAD1D
`define CUBE_LUT_AD21 16'hAD1E
`define CUBE_LUT_AD22 16'hAD1F
`define CUBE_LUT_AD23 16'hAD20
`define CUBE_LUT_AD24 16'hAD21
`define CUBE_LUT_AD25 16'hAD22
`define CUBE_LUT_AD26 16'hAD23
`define CUBE_LUT_AD27 16'hAD24
`define CUBE_LUT_AD28 16'hAD25
`define CUBE_LUT_AD29 16'hAD26
`define CUBE_LUT_AD2A 16'hAD27
`define CUBE_LUT_AD2B 16'hAD28
`define CUBE_LUT_AD2C 16'hAD29
`define CUBE_LUT_AD2D 16'hAD2A
`define CUBE_LUT_AD2E 16'hAD2B
`define CUBE_LUT_AD2F 16'hAD2C
`define CUBE_LUT_AD30 16'hAD2D
`define CUBE_LUT_AD31 16'hAD2E
`define CUBE_LUT_AD32 16'hAD2F
`define CUBE_LUT_AD33 16'hAD30
`define CUBE_LUT_AD34 16'hAD31
`define CUBE_LUT_AD35 16'hAD32
`define CUBE_LUT_AD36 16'hAD33
`define CUBE_LUT_AD37 16'hAD34
`define CUBE_LUT_AD38 16'hAD35
`define CUBE_LUT_AD39 16'hAD36
`define CUBE_LUT_AD3A 16'hAD37
`define CUBE_LUT_AD3B 16'hAD38
`define CUBE_LUT_AD3C 16'hAD39
`define CUBE_LUT_AD3D 16'hAD3A
`define CUBE_LUT_AD3E 16'hAD3B
`define CUBE_LUT_AD3F 16'hAD3C
`define CUBE_LUT_AD40 16'hAD3D
`define CUBE_LUT_AD41 16'hAD3E
`define CUBE_LUT_AD42 16'hAD3F
`define CUBE_LUT_AD43 16'hAD40
`define CUBE_LUT_AD44 16'hAD41
`define CUBE_LUT_AD45 16'hAD42
`define CUBE_LUT_AD46 16'hAD43
`define CUBE_LUT_AD47 16'hAD44
`define CUBE_LUT_AD48 16'hAD45
`define CUBE_LUT_AD49 16'hAD46
`define CUBE_LUT_AD4A 16'hAD47
`define CUBE_LUT_AD4B 16'hAD48
`define CUBE_LUT_AD4C 16'hAD49
`define CUBE_LUT_AD4D 16'hAD4A
`define CUBE_LUT_AD4E 16'hAD4B
`define CUBE_LUT_AD4F 16'hAD4C
`define CUBE_LUT_AD50 16'hAD4D
`define CUBE_LUT_AD51 16'hAD4E
`define CUBE_LUT_AD52 16'hAD4F
`define CUBE_LUT_AD53 16'hAD50
`define CUBE_LUT_AD54 16'hAD51
`define CUBE_LUT_AD55 16'hAD52
`define CUBE_LUT_AD56 16'hAD53
`define CUBE_LUT_AD57 16'hAD54
`define CUBE_LUT_AD58 16'hAD55
`define CUBE_LUT_AD59 16'hAD56
`define CUBE_LUT_AD5A 16'hAD57
`define CUBE_LUT_AD5B 16'hAD58
`define CUBE_LUT_AD5C 16'hAD59
`define CUBE_LUT_AD5D 16'hAD5A
`define CUBE_LUT_AD5E 16'hAD5B
`define CUBE_LUT_AD5F 16'hAD5C
`define CUBE_LUT_AD60 16'hAD5D
`define CUBE_LUT_AD61 16'hAD5E
`define CUBE_LUT_AD62 16'hAD5F
`define CUBE_LUT_AD63 16'hAD60
`define CUBE_LUT_AD64 16'hAD61
`define CUBE_LUT_AD65 16'hAD62
`define CUBE_LUT_AD66 16'hAD63
`define CUBE_LUT_AD67 16'hAD64
`define CUBE_LUT_AD68 16'hAD65
`define CUBE_LUT_AD69 16'hAD66
`define CUBE_LUT_AD6A 16'hAD67
`define CUBE_LUT_AD6B 16'hAD68
`define CUBE_LUT_AD6C 16'hAD69
`define CUBE_LUT_AD6D 16'hAD6A
`define CUBE_LUT_AD6E 16'hAD6B
`define CUBE_LUT_AD6F 16'hAD6C
`define CUBE_LUT_AD70 16'hAD6D
`define CUBE_LUT_AD71 16'hAD6E
`define CUBE_LUT_AD72 16'hAD6F
`define CUBE_LUT_AD73 16'hAD70
`define CUBE_LUT_AD74 16'hAD71
`define CUBE_LUT_AD75 16'hAD72
`define CUBE_LUT_AD76 16'hAD73
`define CUBE_LUT_AD77 16'hAD74
`define CUBE_LUT_AD78 16'hAD75
`define CUBE_LUT_AD79 16'hAD76
`define CUBE_LUT_AD7A 16'hAD77
`define CUBE_LUT_AD7B 16'hAD78
`define CUBE_LUT_AD7C 16'hAD79
`define CUBE_LUT_AD7D 16'hAD7A
`define CUBE_LUT_AD7E 16'hAD7B
`define CUBE_LUT_AD7F 16'hAD7C
`define CUBE_LUT_AD80 16'hAD7D
`define CUBE_LUT_AD81 16'hAD7E
`define CUBE_LUT_AD82 16'hAD7F
`define CUBE_LUT_AD83 16'hAD80
`define CUBE_LUT_AD84 16'hAD81
`define CUBE_LUT_AD85 16'hAD82
`define CUBE_LUT_AD86 16'hAD82
`define CUBE_LUT_AD87 16'hAD83
`define CUBE_LUT_AD88 16'hAD84
`define CUBE_LUT_AD89 16'hAD85
`define CUBE_LUT_AD8A 16'hAD86
`define CUBE_LUT_AD8B 16'hAD87
`define CUBE_LUT_AD8C 16'hAD88
`define CUBE_LUT_AD8D 16'hAD89
`define CUBE_LUT_AD8E 16'hAD8A
`define CUBE_LUT_AD8F 16'hAD8B
`define CUBE_LUT_AD90 16'hAD8C
`define CUBE_LUT_AD91 16'hAD8D
`define CUBE_LUT_AD92 16'hAD8E
`define CUBE_LUT_AD93 16'hAD8F
`define CUBE_LUT_AD94 16'hAD90
`define CUBE_LUT_AD95 16'hAD91
`define CUBE_LUT_AD96 16'hAD92
`define CUBE_LUT_AD97 16'hAD93
`define CUBE_LUT_AD98 16'hAD94
`define CUBE_LUT_AD99 16'hAD95
`define CUBE_LUT_AD9A 16'hAD96
`define CUBE_LUT_AD9B 16'hAD97
`define CUBE_LUT_AD9C 16'hAD98
`define CUBE_LUT_AD9D 16'hAD99
`define CUBE_LUT_AD9E 16'hAD9A
`define CUBE_LUT_AD9F 16'hAD9B
`define CUBE_LUT_ADA0 16'hAD9C
`define CUBE_LUT_ADA1 16'hAD9D
`define CUBE_LUT_ADA2 16'hAD9E
`define CUBE_LUT_ADA3 16'hAD9F
`define CUBE_LUT_ADA4 16'hADA0
`define CUBE_LUT_ADA5 16'hADA1
`define CUBE_LUT_ADA6 16'hADA2
`define CUBE_LUT_ADA7 16'hADA3
`define CUBE_LUT_ADA8 16'hADA4
`define CUBE_LUT_ADA9 16'hADA5
`define CUBE_LUT_ADAA 16'hADA6
`define CUBE_LUT_ADAB 16'hADA7
`define CUBE_LUT_ADAC 16'hADA8
`define CUBE_LUT_ADAD 16'hADA9
`define CUBE_LUT_ADAE 16'hADAA
`define CUBE_LUT_ADAF 16'hADAB
`define CUBE_LUT_ADB0 16'hADAC
`define CUBE_LUT_ADB1 16'hADAD
`define CUBE_LUT_ADB2 16'hADAE
`define CUBE_LUT_ADB3 16'hADAF
`define CUBE_LUT_ADB4 16'hADB0
`define CUBE_LUT_ADB5 16'hADB1
`define CUBE_LUT_ADB6 16'hADB2
`define CUBE_LUT_ADB7 16'hADB3
`define CUBE_LUT_ADB8 16'hADB4
`define CUBE_LUT_ADB9 16'hADB5
`define CUBE_LUT_ADBA 16'hADB6
`define CUBE_LUT_ADBB 16'hADB7
`define CUBE_LUT_ADBC 16'hADB8
`define CUBE_LUT_ADBD 16'hADB9
`define CUBE_LUT_ADBE 16'hADBA
`define CUBE_LUT_ADBF 16'hADBB
`define CUBE_LUT_ADC0 16'hADBC
`define CUBE_LUT_ADC1 16'hADBD
`define CUBE_LUT_ADC2 16'hADBE
`define CUBE_LUT_ADC3 16'hADBF
`define CUBE_LUT_ADC4 16'hADC0
`define CUBE_LUT_ADC5 16'hADC1
`define CUBE_LUT_ADC6 16'hADC2
`define CUBE_LUT_ADC7 16'hADC3
`define CUBE_LUT_ADC8 16'hADC4
`define CUBE_LUT_ADC9 16'hADC5
`define CUBE_LUT_ADCA 16'hADC6
`define CUBE_LUT_ADCB 16'hADC7
`define CUBE_LUT_ADCC 16'hADC8
`define CUBE_LUT_ADCD 16'hADC9
`define CUBE_LUT_ADCE 16'hADCA
`define CUBE_LUT_ADCF 16'hADCB
`define CUBE_LUT_ADD0 16'hADCC
`define CUBE_LUT_ADD1 16'hADCD
`define CUBE_LUT_ADD2 16'hADCE
`define CUBE_LUT_ADD3 16'hADCF
`define CUBE_LUT_ADD4 16'hADD0
`define CUBE_LUT_ADD5 16'hADD1
`define CUBE_LUT_ADD6 16'hADD2
`define CUBE_LUT_ADD7 16'hADD3
`define CUBE_LUT_ADD8 16'hADD4
`define CUBE_LUT_ADD9 16'hADD5
`define CUBE_LUT_ADDA 16'hADD6
`define CUBE_LUT_ADDB 16'hADD7
`define CUBE_LUT_ADDC 16'hADD8
`define CUBE_LUT_ADDD 16'hADD9
`define CUBE_LUT_ADDE 16'hADDA
`define CUBE_LUT_ADDF 16'hADDB
`define CUBE_LUT_ADE0 16'hADDC
`define CUBE_LUT_ADE1 16'hADDD
`define CUBE_LUT_ADE2 16'hADDE
`define CUBE_LUT_ADE3 16'hADDF
`define CUBE_LUT_ADE4 16'hADE0
`define CUBE_LUT_ADE5 16'hADE1
`define CUBE_LUT_ADE6 16'hADE2
`define CUBE_LUT_ADE7 16'hADE3
`define CUBE_LUT_ADE8 16'hADE4
`define CUBE_LUT_ADE9 16'hADE5
`define CUBE_LUT_ADEA 16'hADE6
`define CUBE_LUT_ADEB 16'hADE7
`define CUBE_LUT_ADEC 16'hADE8
`define CUBE_LUT_ADED 16'hADE9
`define CUBE_LUT_ADEE 16'hADEA
`define CUBE_LUT_ADEF 16'hADEB
`define CUBE_LUT_ADF0 16'hADEC
`define CUBE_LUT_ADF1 16'hADED
`define CUBE_LUT_ADF2 16'hADEE
`define CUBE_LUT_ADF3 16'hADEF
`define CUBE_LUT_ADF4 16'hADF0
`define CUBE_LUT_ADF5 16'hADF1
`define CUBE_LUT_ADF6 16'hADF2
`define CUBE_LUT_ADF7 16'hADF3
`define CUBE_LUT_ADF8 16'hADF4
`define CUBE_LUT_ADF9 16'hADF5
`define CUBE_LUT_ADFA 16'hADF6
`define CUBE_LUT_ADFB 16'hADF7
`define CUBE_LUT_ADFC 16'hADF8
`define CUBE_LUT_ADFD 16'hADF9
`define CUBE_LUT_ADFE 16'hADFA
`define CUBE_LUT_ADFF 16'hADFB
`define CUBE_LUT_AE00 16'hADFC
`define CUBE_LUT_AE01 16'hADFD
`define CUBE_LUT_AE02 16'hADFD
`define CUBE_LUT_AE03 16'hADFE
`define CUBE_LUT_AE04 16'hADFF
`define CUBE_LUT_AE05 16'hAE00
`define CUBE_LUT_AE06 16'hAE01
`define CUBE_LUT_AE07 16'hAE02
`define CUBE_LUT_AE08 16'hAE03
`define CUBE_LUT_AE09 16'hAE04
`define CUBE_LUT_AE0A 16'hAE05
`define CUBE_LUT_AE0B 16'hAE06
`define CUBE_LUT_AE0C 16'hAE07
`define CUBE_LUT_AE0D 16'hAE08
`define CUBE_LUT_AE0E 16'hAE09
`define CUBE_LUT_AE0F 16'hAE0A
`define CUBE_LUT_AE10 16'hAE0B
`define CUBE_LUT_AE11 16'hAE0C
`define CUBE_LUT_AE12 16'hAE0D
`define CUBE_LUT_AE13 16'hAE0E
`define CUBE_LUT_AE14 16'hAE0F
`define CUBE_LUT_AE15 16'hAE10
`define CUBE_LUT_AE16 16'hAE11
`define CUBE_LUT_AE17 16'hAE12
`define CUBE_LUT_AE18 16'hAE13
`define CUBE_LUT_AE19 16'hAE14
`define CUBE_LUT_AE1A 16'hAE15
`define CUBE_LUT_AE1B 16'hAE16
`define CUBE_LUT_AE1C 16'hAE17
`define CUBE_LUT_AE1D 16'hAE18
`define CUBE_LUT_AE1E 16'hAE19
`define CUBE_LUT_AE1F 16'hAE1A
`define CUBE_LUT_AE20 16'hAE1B
`define CUBE_LUT_AE21 16'hAE1C
`define CUBE_LUT_AE22 16'hAE1D
`define CUBE_LUT_AE23 16'hAE1E
`define CUBE_LUT_AE24 16'hAE1F
`define CUBE_LUT_AE25 16'hAE20
`define CUBE_LUT_AE26 16'hAE21
`define CUBE_LUT_AE27 16'hAE22
`define CUBE_LUT_AE28 16'hAE23
`define CUBE_LUT_AE29 16'hAE24
`define CUBE_LUT_AE2A 16'hAE25
`define CUBE_LUT_AE2B 16'hAE26
`define CUBE_LUT_AE2C 16'hAE27
`define CUBE_LUT_AE2D 16'hAE28
`define CUBE_LUT_AE2E 16'hAE29
`define CUBE_LUT_AE2F 16'hAE2A
`define CUBE_LUT_AE30 16'hAE2B
`define CUBE_LUT_AE31 16'hAE2C
`define CUBE_LUT_AE32 16'hAE2D
`define CUBE_LUT_AE33 16'hAE2E
`define CUBE_LUT_AE34 16'hAE2F
`define CUBE_LUT_AE35 16'hAE30
`define CUBE_LUT_AE36 16'hAE31
`define CUBE_LUT_AE37 16'hAE32
`define CUBE_LUT_AE38 16'hAE33
`define CUBE_LUT_AE39 16'hAE34
`define CUBE_LUT_AE3A 16'hAE35
`define CUBE_LUT_AE3B 16'hAE36
`define CUBE_LUT_AE3C 16'hAE37
`define CUBE_LUT_AE3D 16'hAE38
`define CUBE_LUT_AE3E 16'hAE39
`define CUBE_LUT_AE3F 16'hAE3A
`define CUBE_LUT_AE40 16'hAE3B
`define CUBE_LUT_AE41 16'hAE3C
`define CUBE_LUT_AE42 16'hAE3D
`define CUBE_LUT_AE43 16'hAE3E
`define CUBE_LUT_AE44 16'hAE3F
`define CUBE_LUT_AE45 16'hAE40
`define CUBE_LUT_AE46 16'hAE41
`define CUBE_LUT_AE47 16'hAE42
`define CUBE_LUT_AE48 16'hAE43
`define CUBE_LUT_AE49 16'hAE44
`define CUBE_LUT_AE4A 16'hAE45
`define CUBE_LUT_AE4B 16'hAE46
`define CUBE_LUT_AE4C 16'hAE47
`define CUBE_LUT_AE4D 16'hAE48
`define CUBE_LUT_AE4E 16'hAE49
`define CUBE_LUT_AE4F 16'hAE4A
`define CUBE_LUT_AE50 16'hAE4B
`define CUBE_LUT_AE51 16'hAE4C
`define CUBE_LUT_AE52 16'hAE4D
`define CUBE_LUT_AE53 16'hAE4E
`define CUBE_LUT_AE54 16'hAE4F
`define CUBE_LUT_AE55 16'hAE50
`define CUBE_LUT_AE56 16'hAE51
`define CUBE_LUT_AE57 16'hAE52
`define CUBE_LUT_AE58 16'hAE53
`define CUBE_LUT_AE59 16'hAE54
`define CUBE_LUT_AE5A 16'hAE55
`define CUBE_LUT_AE5B 16'hAE56
`define CUBE_LUT_AE5C 16'hAE57
`define CUBE_LUT_AE5D 16'hAE58
`define CUBE_LUT_AE5E 16'hAE59
`define CUBE_LUT_AE5F 16'hAE5A
`define CUBE_LUT_AE60 16'hAE5B
`define CUBE_LUT_AE61 16'hAE5C
`define CUBE_LUT_AE62 16'hAE5D
`define CUBE_LUT_AE63 16'hAE5E
`define CUBE_LUT_AE64 16'hAE5F
`define CUBE_LUT_AE65 16'hAE60
`define CUBE_LUT_AE66 16'hAE61
`define CUBE_LUT_AE67 16'hAE62
`define CUBE_LUT_AE68 16'hAE63
`define CUBE_LUT_AE69 16'hAE64
`define CUBE_LUT_AE6A 16'hAE65
`define CUBE_LUT_AE6B 16'hAE66
`define CUBE_LUT_AE6C 16'hAE67
`define CUBE_LUT_AE6D 16'hAE67
`define CUBE_LUT_AE6E 16'hAE68
`define CUBE_LUT_AE6F 16'hAE69
`define CUBE_LUT_AE70 16'hAE6A
`define CUBE_LUT_AE71 16'hAE6B
`define CUBE_LUT_AE72 16'hAE6C
`define CUBE_LUT_AE73 16'hAE6D
`define CUBE_LUT_AE74 16'hAE6E
`define CUBE_LUT_AE75 16'hAE6F
`define CUBE_LUT_AE76 16'hAE70
`define CUBE_LUT_AE77 16'hAE71
`define CUBE_LUT_AE78 16'hAE72
`define CUBE_LUT_AE79 16'hAE73
`define CUBE_LUT_AE7A 16'hAE74
`define CUBE_LUT_AE7B 16'hAE75
`define CUBE_LUT_AE7C 16'hAE76
`define CUBE_LUT_AE7D 16'hAE77
`define CUBE_LUT_AE7E 16'hAE78
`define CUBE_LUT_AE7F 16'hAE79
`define CUBE_LUT_AE80 16'hAE7A
`define CUBE_LUT_AE81 16'hAE7B
`define CUBE_LUT_AE82 16'hAE7C
`define CUBE_LUT_AE83 16'hAE7D
`define CUBE_LUT_AE84 16'hAE7E
`define CUBE_LUT_AE85 16'hAE7F
`define CUBE_LUT_AE86 16'hAE80
`define CUBE_LUT_AE87 16'hAE81
`define CUBE_LUT_AE88 16'hAE82
`define CUBE_LUT_AE89 16'hAE83
`define CUBE_LUT_AE8A 16'hAE84
`define CUBE_LUT_AE8B 16'hAE85
`define CUBE_LUT_AE8C 16'hAE86
`define CUBE_LUT_AE8D 16'hAE87
`define CUBE_LUT_AE8E 16'hAE88
`define CUBE_LUT_AE8F 16'hAE89
`define CUBE_LUT_AE90 16'hAE8A
`define CUBE_LUT_AE91 16'hAE8B
`define CUBE_LUT_AE92 16'hAE8C
`define CUBE_LUT_AE93 16'hAE8D
`define CUBE_LUT_AE94 16'hAE8E
`define CUBE_LUT_AE95 16'hAE8F
`define CUBE_LUT_AE96 16'hAE90
`define CUBE_LUT_AE97 16'hAE91
`define CUBE_LUT_AE98 16'hAE92
`define CUBE_LUT_AE99 16'hAE93
`define CUBE_LUT_AE9A 16'hAE94
`define CUBE_LUT_AE9B 16'hAE95
`define CUBE_LUT_AE9C 16'hAE96
`define CUBE_LUT_AE9D 16'hAE97
`define CUBE_LUT_AE9E 16'hAE98
`define CUBE_LUT_AE9F 16'hAE99
`define CUBE_LUT_AEA0 16'hAE9A
`define CUBE_LUT_AEA1 16'hAE9B
`define CUBE_LUT_AEA2 16'hAE9C
`define CUBE_LUT_AEA3 16'hAE9D
`define CUBE_LUT_AEA4 16'hAE9E
`define CUBE_LUT_AEA5 16'hAE9F
`define CUBE_LUT_AEA6 16'hAEA0
`define CUBE_LUT_AEA7 16'hAEA1
`define CUBE_LUT_AEA8 16'hAEA2
`define CUBE_LUT_AEA9 16'hAEA3
`define CUBE_LUT_AEAA 16'hAEA4
`define CUBE_LUT_AEAB 16'hAEA5
`define CUBE_LUT_AEAC 16'hAEA6
`define CUBE_LUT_AEAD 16'hAEA7
`define CUBE_LUT_AEAE 16'hAEA8
`define CUBE_LUT_AEAF 16'hAEA9
`define CUBE_LUT_AEB0 16'hAEAA
`define CUBE_LUT_AEB1 16'hAEAB
`define CUBE_LUT_AEB2 16'hAEAC
`define CUBE_LUT_AEB3 16'hAEAD
`define CUBE_LUT_AEB4 16'hAEAE
`define CUBE_LUT_AEB5 16'hAEAF
`define CUBE_LUT_AEB6 16'hAEB0
`define CUBE_LUT_AEB7 16'hAEB1
`define CUBE_LUT_AEB8 16'hAEB2
`define CUBE_LUT_AEB9 16'hAEB3
`define CUBE_LUT_AEBA 16'hAEB4
`define CUBE_LUT_AEBB 16'hAEB5
`define CUBE_LUT_AEBC 16'hAEB6
`define CUBE_LUT_AEBD 16'hAEB7
`define CUBE_LUT_AEBE 16'hAEB8
`define CUBE_LUT_AEBF 16'hAEB9
`define CUBE_LUT_AEC0 16'hAEBA
`define CUBE_LUT_AEC1 16'hAEBB
`define CUBE_LUT_AEC2 16'hAEBC
`define CUBE_LUT_AEC3 16'hAEBD
`define CUBE_LUT_AEC4 16'hAEBE
`define CUBE_LUT_AEC5 16'hAEBF
`define CUBE_LUT_AEC6 16'hAEC0
`define CUBE_LUT_AEC7 16'hAEC1
`define CUBE_LUT_AEC8 16'hAEC2
`define CUBE_LUT_AEC9 16'hAEC3
`define CUBE_LUT_AECA 16'hAEC4
`define CUBE_LUT_AECB 16'hAEC4
`define CUBE_LUT_AECC 16'hAEC5
`define CUBE_LUT_AECD 16'hAEC6
`define CUBE_LUT_AECE 16'hAEC7
`define CUBE_LUT_AECF 16'hAEC8
`define CUBE_LUT_AED0 16'hAEC9
`define CUBE_LUT_AED1 16'hAECA
`define CUBE_LUT_AED2 16'hAECB
`define CUBE_LUT_AED3 16'hAECC
`define CUBE_LUT_AED4 16'hAECD
`define CUBE_LUT_AED5 16'hAECE
`define CUBE_LUT_AED6 16'hAECF
`define CUBE_LUT_AED7 16'hAED0
`define CUBE_LUT_AED8 16'hAED1
`define CUBE_LUT_AED9 16'hAED2
`define CUBE_LUT_AEDA 16'hAED3
`define CUBE_LUT_AEDB 16'hAED4
`define CUBE_LUT_AEDC 16'hAED5
`define CUBE_LUT_AEDD 16'hAED6
`define CUBE_LUT_AEDE 16'hAED7
`define CUBE_LUT_AEDF 16'hAED8
`define CUBE_LUT_AEE0 16'hAED9
`define CUBE_LUT_AEE1 16'hAEDA
`define CUBE_LUT_AEE2 16'hAEDB
`define CUBE_LUT_AEE3 16'hAEDC
`define CUBE_LUT_AEE4 16'hAEDD
`define CUBE_LUT_AEE5 16'hAEDE
`define CUBE_LUT_AEE6 16'hAEDF
`define CUBE_LUT_AEE7 16'hAEE0
`define CUBE_LUT_AEE8 16'hAEE1
`define CUBE_LUT_AEE9 16'hAEE2
`define CUBE_LUT_AEEA 16'hAEE3
`define CUBE_LUT_AEEB 16'hAEE4
`define CUBE_LUT_AEEC 16'hAEE5
`define CUBE_LUT_AEED 16'hAEE6
`define CUBE_LUT_AEEE 16'hAEE7
`define CUBE_LUT_AEEF 16'hAEE8
`define CUBE_LUT_AEF0 16'hAEE9
`define CUBE_LUT_AEF1 16'hAEEA
`define CUBE_LUT_AEF2 16'hAEEB
`define CUBE_LUT_AEF3 16'hAEEC
`define CUBE_LUT_AEF4 16'hAEED
`define CUBE_LUT_AEF5 16'hAEEE
`define CUBE_LUT_AEF6 16'hAEEF
`define CUBE_LUT_AEF7 16'hAEF0
`define CUBE_LUT_AEF8 16'hAEF1
`define CUBE_LUT_AEF9 16'hAEF2
`define CUBE_LUT_AEFA 16'hAEF3
`define CUBE_LUT_AEFB 16'hAEF4
`define CUBE_LUT_AEFC 16'hAEF5
`define CUBE_LUT_AEFD 16'hAEF6
`define CUBE_LUT_AEFE 16'hAEF7
`define CUBE_LUT_AEFF 16'hAEF8
`define CUBE_LUT_AF00 16'hAEF9
`define CUBE_LUT_AF01 16'hAEFA
`define CUBE_LUT_AF02 16'hAEFB
`define CUBE_LUT_AF03 16'hAEFC
`define CUBE_LUT_AF04 16'hAEFD
`define CUBE_LUT_AF05 16'hAEFE
`define CUBE_LUT_AF06 16'hAEFF
`define CUBE_LUT_AF07 16'hAF00
`define CUBE_LUT_AF08 16'hAF01
`define CUBE_LUT_AF09 16'hAF02
`define CUBE_LUT_AF0A 16'hAF03
`define CUBE_LUT_AF0B 16'hAF04
`define CUBE_LUT_AF0C 16'hAF05
`define CUBE_LUT_AF0D 16'hAF06
`define CUBE_LUT_AF0E 16'hAF07
`define CUBE_LUT_AF0F 16'hAF08
`define CUBE_LUT_AF10 16'hAF09
`define CUBE_LUT_AF11 16'hAF0A
`define CUBE_LUT_AF12 16'hAF0B
`define CUBE_LUT_AF13 16'hAF0C
`define CUBE_LUT_AF14 16'hAF0D
`define CUBE_LUT_AF15 16'hAF0E
`define CUBE_LUT_AF16 16'hAF0F
`define CUBE_LUT_AF17 16'hAF10
`define CUBE_LUT_AF18 16'hAF11
`define CUBE_LUT_AF19 16'hAF12
`define CUBE_LUT_AF1A 16'hAF13
`define CUBE_LUT_AF1B 16'hAF14
`define CUBE_LUT_AF1C 16'hAF15
`define CUBE_LUT_AF1D 16'hAF16
`define CUBE_LUT_AF1E 16'hAF17
`define CUBE_LUT_AF1F 16'hAF18
`define CUBE_LUT_AF20 16'hAF19
`define CUBE_LUT_AF21 16'hAF19
`define CUBE_LUT_AF22 16'hAF1A
`define CUBE_LUT_AF23 16'hAF1B
`define CUBE_LUT_AF24 16'hAF1C
`define CUBE_LUT_AF25 16'hAF1D
`define CUBE_LUT_AF26 16'hAF1E
`define CUBE_LUT_AF27 16'hAF1F
`define CUBE_LUT_AF28 16'hAF20
`define CUBE_LUT_AF29 16'hAF21
`define CUBE_LUT_AF2A 16'hAF22
`define CUBE_LUT_AF2B 16'hAF23
`define CUBE_LUT_AF2C 16'hAF24
`define CUBE_LUT_AF2D 16'hAF25
`define CUBE_LUT_AF2E 16'hAF26
`define CUBE_LUT_AF2F 16'hAF27
`define CUBE_LUT_AF30 16'hAF28
`define CUBE_LUT_AF31 16'hAF29
`define CUBE_LUT_AF32 16'hAF2A
`define CUBE_LUT_AF33 16'hAF2B
`define CUBE_LUT_AF34 16'hAF2C
`define CUBE_LUT_AF35 16'hAF2D
`define CUBE_LUT_AF36 16'hAF2E
`define CUBE_LUT_AF37 16'hAF2F
`define CUBE_LUT_AF38 16'hAF30
`define CUBE_LUT_AF39 16'hAF31
`define CUBE_LUT_AF3A 16'hAF32
`define CUBE_LUT_AF3B 16'hAF33
`define CUBE_LUT_AF3C 16'hAF34
`define CUBE_LUT_AF3D 16'hAF35
`define CUBE_LUT_AF3E 16'hAF36
`define CUBE_LUT_AF3F 16'hAF37
`define CUBE_LUT_AF40 16'hAF38
`define CUBE_LUT_AF41 16'hAF39
`define CUBE_LUT_AF42 16'hAF3A
`define CUBE_LUT_AF43 16'hAF3B
`define CUBE_LUT_AF44 16'hAF3C
`define CUBE_LUT_AF45 16'hAF3D
`define CUBE_LUT_AF46 16'hAF3E
`define CUBE_LUT_AF47 16'hAF3F
`define CUBE_LUT_AF48 16'hAF40
`define CUBE_LUT_AF49 16'hAF41
`define CUBE_LUT_AF4A 16'hAF42
`define CUBE_LUT_AF4B 16'hAF43
`define CUBE_LUT_AF4C 16'hAF44
`define CUBE_LUT_AF4D 16'hAF45
`define CUBE_LUT_AF4E 16'hAF46
`define CUBE_LUT_AF4F 16'hAF47
`define CUBE_LUT_AF50 16'hAF48
`define CUBE_LUT_AF51 16'hAF49
`define CUBE_LUT_AF52 16'hAF4A
`define CUBE_LUT_AF53 16'hAF4B
`define CUBE_LUT_AF54 16'hAF4C
`define CUBE_LUT_AF55 16'hAF4D
`define CUBE_LUT_AF56 16'hAF4E
`define CUBE_LUT_AF57 16'hAF4F
`define CUBE_LUT_AF58 16'hAF50
`define CUBE_LUT_AF59 16'hAF51
`define CUBE_LUT_AF5A 16'hAF52
`define CUBE_LUT_AF5B 16'hAF53
`define CUBE_LUT_AF5C 16'hAF54
`define CUBE_LUT_AF5D 16'hAF55
`define CUBE_LUT_AF5E 16'hAF56
`define CUBE_LUT_AF5F 16'hAF57
`define CUBE_LUT_AF60 16'hAF58
`define CUBE_LUT_AF61 16'hAF59
`define CUBE_LUT_AF62 16'hAF5A
`define CUBE_LUT_AF63 16'hAF5B
`define CUBE_LUT_AF64 16'hAF5C
`define CUBE_LUT_AF65 16'hAF5D
`define CUBE_LUT_AF66 16'hAF5E
`define CUBE_LUT_AF67 16'hAF5F
`define CUBE_LUT_AF68 16'hAF60
`define CUBE_LUT_AF69 16'hAF61
`define CUBE_LUT_AF6A 16'hAF62
`define CUBE_LUT_AF6B 16'hAF63
`define CUBE_LUT_AF6C 16'hAF64
`define CUBE_LUT_AF6D 16'hAF65
`define CUBE_LUT_AF6E 16'hAF66
`define CUBE_LUT_AF6F 16'hAF66
`define CUBE_LUT_AF70 16'hAF67
`define CUBE_LUT_AF71 16'hAF68
`define CUBE_LUT_AF72 16'hAF69
`define CUBE_LUT_AF73 16'hAF6A
`define CUBE_LUT_AF74 16'hAF6B
`define CUBE_LUT_AF75 16'hAF6C
`define CUBE_LUT_AF76 16'hAF6D
`define CUBE_LUT_AF77 16'hAF6E
`define CUBE_LUT_AF78 16'hAF6F
`define CUBE_LUT_AF79 16'hAF70
`define CUBE_LUT_AF7A 16'hAF71
`define CUBE_LUT_AF7B 16'hAF72
`define CUBE_LUT_AF7C 16'hAF73
`define CUBE_LUT_AF7D 16'hAF74
`define CUBE_LUT_AF7E 16'hAF75
`define CUBE_LUT_AF7F 16'hAF76
`define CUBE_LUT_AF80 16'hAF77
`define CUBE_LUT_AF81 16'hAF78
`define CUBE_LUT_AF82 16'hAF79
`define CUBE_LUT_AF83 16'hAF7A
`define CUBE_LUT_AF84 16'hAF7B
`define CUBE_LUT_AF85 16'hAF7C
`define CUBE_LUT_AF86 16'hAF7D
`define CUBE_LUT_AF87 16'hAF7E
`define CUBE_LUT_AF88 16'hAF7F
`define CUBE_LUT_AF89 16'hAF80
`define CUBE_LUT_AF8A 16'hAF81
`define CUBE_LUT_AF8B 16'hAF82
`define CUBE_LUT_AF8C 16'hAF83
`define CUBE_LUT_AF8D 16'hAF84
`define CUBE_LUT_AF8E 16'hAF85
`define CUBE_LUT_AF8F 16'hAF86
`define CUBE_LUT_AF90 16'hAF87
`define CUBE_LUT_AF91 16'hAF88
`define CUBE_LUT_AF92 16'hAF89
`define CUBE_LUT_AF93 16'hAF8A
`define CUBE_LUT_AF94 16'hAF8B
`define CUBE_LUT_AF95 16'hAF8C
`define CUBE_LUT_AF96 16'hAF8D
`define CUBE_LUT_AF97 16'hAF8E
`define CUBE_LUT_AF98 16'hAF8F
`define CUBE_LUT_AF99 16'hAF90
`define CUBE_LUT_AF9A 16'hAF91
`define CUBE_LUT_AF9B 16'hAF92
`define CUBE_LUT_AF9C 16'hAF93
`define CUBE_LUT_AF9D 16'hAF94
`define CUBE_LUT_AF9E 16'hAF95
`define CUBE_LUT_AF9F 16'hAF96
`define CUBE_LUT_AFA0 16'hAF97
`define CUBE_LUT_AFA1 16'hAF98
`define CUBE_LUT_AFA2 16'hAF99
`define CUBE_LUT_AFA3 16'hAF9A
`define CUBE_LUT_AFA4 16'hAF9B
`define CUBE_LUT_AFA5 16'hAF9C
`define CUBE_LUT_AFA6 16'hAF9D
`define CUBE_LUT_AFA7 16'hAF9E
`define CUBE_LUT_AFA8 16'hAF9F
`define CUBE_LUT_AFA9 16'hAFA0
`define CUBE_LUT_AFAA 16'hAFA1
`define CUBE_LUT_AFAB 16'hAFA2
`define CUBE_LUT_AFAC 16'hAFA3
`define CUBE_LUT_AFAD 16'hAFA4
`define CUBE_LUT_AFAE 16'hAFA5
`define CUBE_LUT_AFAF 16'hAFA6
`define CUBE_LUT_AFB0 16'hAFA7
`define CUBE_LUT_AFB1 16'hAFA8
`define CUBE_LUT_AFB2 16'hAFA9
`define CUBE_LUT_AFB3 16'hAFAA
`define CUBE_LUT_AFB4 16'hAFAB
`define CUBE_LUT_AFB5 16'hAFAC
`define CUBE_LUT_AFB6 16'hAFAD
`define CUBE_LUT_AFB7 16'hAFAD
`define CUBE_LUT_AFB8 16'hAFAE
`define CUBE_LUT_AFB9 16'hAFAF
`define CUBE_LUT_AFBA 16'hAFB0
`define CUBE_LUT_AFBB 16'hAFB1
`define CUBE_LUT_AFBC 16'hAFB2
`define CUBE_LUT_AFBD 16'hAFB3
`define CUBE_LUT_AFBE 16'hAFB4
`define CUBE_LUT_AFBF 16'hAFB5
`define CUBE_LUT_AFC0 16'hAFB6
`define CUBE_LUT_AFC1 16'hAFB7
`define CUBE_LUT_AFC2 16'hAFB8
`define CUBE_LUT_AFC3 16'hAFB9
`define CUBE_LUT_AFC4 16'hAFBA
`define CUBE_LUT_AFC5 16'hAFBB
`define CUBE_LUT_AFC6 16'hAFBC
`define CUBE_LUT_AFC7 16'hAFBD
`define CUBE_LUT_AFC8 16'hAFBE
`define CUBE_LUT_AFC9 16'hAFBF
`define CUBE_LUT_AFCA 16'hAFC0
`define CUBE_LUT_AFCB 16'hAFC1
`define CUBE_LUT_AFCC 16'hAFC2
`define CUBE_LUT_AFCD 16'hAFC3
`define CUBE_LUT_AFCE 16'hAFC4
`define CUBE_LUT_AFCF 16'hAFC5
`define CUBE_LUT_AFD0 16'hAFC6
`define CUBE_LUT_AFD1 16'hAFC7
`define CUBE_LUT_AFD2 16'hAFC8
`define CUBE_LUT_AFD3 16'hAFC9
`define CUBE_LUT_AFD4 16'hAFCA
`define CUBE_LUT_AFD5 16'hAFCB
`define CUBE_LUT_AFD6 16'hAFCC
`define CUBE_LUT_AFD7 16'hAFCD
`define CUBE_LUT_AFD8 16'hAFCE
`define CUBE_LUT_AFD9 16'hAFCF
`define CUBE_LUT_AFDA 16'hAFD0
`define CUBE_LUT_AFDB 16'hAFD1
`define CUBE_LUT_AFDC 16'hAFD2
`define CUBE_LUT_AFDD 16'hAFD3
`define CUBE_LUT_AFDE 16'hAFD4
`define CUBE_LUT_AFDF 16'hAFD5
`define CUBE_LUT_AFE0 16'hAFD6
`define CUBE_LUT_AFE1 16'hAFD7
`define CUBE_LUT_AFE2 16'hAFD8
`define CUBE_LUT_AFE3 16'hAFD9
`define CUBE_LUT_AFE4 16'hAFDA
`define CUBE_LUT_AFE5 16'hAFDB
`define CUBE_LUT_AFE6 16'hAFDC
`define CUBE_LUT_AFE7 16'hAFDD
`define CUBE_LUT_AFE8 16'hAFDE
`define CUBE_LUT_AFE9 16'hAFDF
`define CUBE_LUT_AFEA 16'hAFE0
`define CUBE_LUT_AFEB 16'hAFE1
`define CUBE_LUT_AFEC 16'hAFE2
`define CUBE_LUT_AFED 16'hAFE3
`define CUBE_LUT_AFEE 16'hAFE4
`define CUBE_LUT_AFEF 16'hAFE5
`define CUBE_LUT_AFF0 16'hAFE6
`define CUBE_LUT_AFF1 16'hAFE7
`define CUBE_LUT_AFF2 16'hAFE8
`define CUBE_LUT_AFF3 16'hAFE9
`define CUBE_LUT_AFF4 16'hAFEA
`define CUBE_LUT_AFF5 16'hAFEB
`define CUBE_LUT_AFF6 16'hAFEC
`define CUBE_LUT_AFF7 16'hAFED
`define CUBE_LUT_AFF8 16'hAFEE
`define CUBE_LUT_AFF9 16'hAFEF
`define CUBE_LUT_AFFA 16'hAFEF
`define CUBE_LUT_AFFB 16'hAFF0
`define CUBE_LUT_AFFC 16'hAFF1
`define CUBE_LUT_AFFD 16'hAFF2
`define CUBE_LUT_AFFE 16'hAFF3
`define CUBE_LUT_AFFF 16'hAFF4
`define CUBE_LUT_B000 16'hAFF5
`define CUBE_LUT_B001 16'hAFF7
`define CUBE_LUT_B002 16'hAFF9
`define CUBE_LUT_B003 16'hAFFB
`define CUBE_LUT_B004 16'hAFFD
`define CUBE_LUT_B005 16'hAFFF
`define CUBE_LUT_B006 16'hB001
`define CUBE_LUT_B007 16'hB002
`define CUBE_LUT_B008 16'hB003
`define CUBE_LUT_B009 16'hB004
`define CUBE_LUT_B00A 16'hB005
`define CUBE_LUT_B00B 16'hB006
`define CUBE_LUT_B00C 16'hB007
`define CUBE_LUT_B00D 16'hB007
`define CUBE_LUT_B00E 16'hB008
`define CUBE_LUT_B00F 16'hB009
`define CUBE_LUT_B010 16'hB00A
`define CUBE_LUT_B011 16'hB00B
`define CUBE_LUT_B012 16'hB00C
`define CUBE_LUT_B013 16'hB00D
`define CUBE_LUT_B014 16'hB00E
`define CUBE_LUT_B015 16'hB00F
`define CUBE_LUT_B016 16'hB010
`define CUBE_LUT_B017 16'hB011
`define CUBE_LUT_B018 16'hB012
`define CUBE_LUT_B019 16'hB013
`define CUBE_LUT_B01A 16'hB014
`define CUBE_LUT_B01B 16'hB015
`define CUBE_LUT_B01C 16'hB016
`define CUBE_LUT_B01D 16'hB017
`define CUBE_LUT_B01E 16'hB018
`define CUBE_LUT_B01F 16'hB019
`define CUBE_LUT_B020 16'hB01A
`define CUBE_LUT_B021 16'hB01B
`define CUBE_LUT_B022 16'hB01C
`define CUBE_LUT_B023 16'hB01D
`define CUBE_LUT_B024 16'hB01E
`define CUBE_LUT_B025 16'hB01F
`define CUBE_LUT_B026 16'hB020
`define CUBE_LUT_B027 16'hB021
`define CUBE_LUT_B028 16'hB022
`define CUBE_LUT_B029 16'hB023
`define CUBE_LUT_B02A 16'hB024
`define CUBE_LUT_B02B 16'hB025
`define CUBE_LUT_B02C 16'hB026
`define CUBE_LUT_B02D 16'hB027
`define CUBE_LUT_B02E 16'hB028
`define CUBE_LUT_B02F 16'hB029
`define CUBE_LUT_B030 16'hB02A
`define CUBE_LUT_B031 16'hB02B
`define CUBE_LUT_B032 16'hB02C
`define CUBE_LUT_B033 16'hB02D
`define CUBE_LUT_B034 16'hB02E
`define CUBE_LUT_B035 16'hB02F
`define CUBE_LUT_B036 16'hB030
`define CUBE_LUT_B037 16'hB031
`define CUBE_LUT_B038 16'hB032
`define CUBE_LUT_B039 16'hB033
`define CUBE_LUT_B03A 16'hB034
`define CUBE_LUT_B03B 16'hB035
`define CUBE_LUT_B03C 16'hB036
`define CUBE_LUT_B03D 16'hB037
`define CUBE_LUT_B03E 16'hB038
`define CUBE_LUT_B03F 16'hB039
`define CUBE_LUT_B040 16'hB03A
`define CUBE_LUT_B041 16'hB03B
`define CUBE_LUT_B042 16'hB03C
`define CUBE_LUT_B043 16'hB03D
`define CUBE_LUT_B044 16'hB03E
`define CUBE_LUT_B045 16'hB03F
`define CUBE_LUT_B046 16'hB040
`define CUBE_LUT_B047 16'hB041
`define CUBE_LUT_B048 16'hB042
`define CUBE_LUT_B049 16'hB042
`define CUBE_LUT_B04A 16'hB043
`define CUBE_LUT_B04B 16'hB044
`define CUBE_LUT_B04C 16'hB045
`define CUBE_LUT_B04D 16'hB046
`define CUBE_LUT_B04E 16'hB047
`define CUBE_LUT_B04F 16'hB048
`define CUBE_LUT_B050 16'hB049
`define CUBE_LUT_B051 16'hB04A
`define CUBE_LUT_B052 16'hB04B
`define CUBE_LUT_B053 16'hB04C
`define CUBE_LUT_B054 16'hB04D
`define CUBE_LUT_B055 16'hB04E
`define CUBE_LUT_B056 16'hB04F
`define CUBE_LUT_B057 16'hB050
`define CUBE_LUT_B058 16'hB051
`define CUBE_LUT_B059 16'hB052
`define CUBE_LUT_B05A 16'hB053
`define CUBE_LUT_B05B 16'hB054
`define CUBE_LUT_B05C 16'hB055
`define CUBE_LUT_B05D 16'hB056
`define CUBE_LUT_B05E 16'hB057
`define CUBE_LUT_B05F 16'hB058
`define CUBE_LUT_B060 16'hB059
`define CUBE_LUT_B061 16'hB05A
`define CUBE_LUT_B062 16'hB05B
`define CUBE_LUT_B063 16'hB05C
`define CUBE_LUT_B064 16'hB05D
`define CUBE_LUT_B065 16'hB05E
`define CUBE_LUT_B066 16'hB05F
`define CUBE_LUT_B067 16'hB060
`define CUBE_LUT_B068 16'hB061
`define CUBE_LUT_B069 16'hB062
`define CUBE_LUT_B06A 16'hB063
`define CUBE_LUT_B06B 16'hB064
`define CUBE_LUT_B06C 16'hB065
`define CUBE_LUT_B06D 16'hB066
`define CUBE_LUT_B06E 16'hB067
`define CUBE_LUT_B06F 16'hB068
`define CUBE_LUT_B070 16'hB069
`define CUBE_LUT_B071 16'hB06A
`define CUBE_LUT_B072 16'hB06B
`define CUBE_LUT_B073 16'hB06C
`define CUBE_LUT_B074 16'hB06D
`define CUBE_LUT_B075 16'hB06E
`define CUBE_LUT_B076 16'hB06F
`define CUBE_LUT_B077 16'hB070
`define CUBE_LUT_B078 16'hB071
`define CUBE_LUT_B079 16'hB072
`define CUBE_LUT_B07A 16'hB073
`define CUBE_LUT_B07B 16'hB074
`define CUBE_LUT_B07C 16'hB075
`define CUBE_LUT_B07D 16'hB076
`define CUBE_LUT_B07E 16'hB077
`define CUBE_LUT_B07F 16'hB077
`define CUBE_LUT_B080 16'hB078
`define CUBE_LUT_B081 16'hB079
`define CUBE_LUT_B082 16'hB07A
`define CUBE_LUT_B083 16'hB07B
`define CUBE_LUT_B084 16'hB07C
`define CUBE_LUT_B085 16'hB07D
`define CUBE_LUT_B086 16'hB07E
`define CUBE_LUT_B087 16'hB07F
`define CUBE_LUT_B088 16'hB080
`define CUBE_LUT_B089 16'hB081
`define CUBE_LUT_B08A 16'hB082
`define CUBE_LUT_B08B 16'hB083
`define CUBE_LUT_B08C 16'hB084
`define CUBE_LUT_B08D 16'hB085
`define CUBE_LUT_B08E 16'hB086
`define CUBE_LUT_B08F 16'hB087
`define CUBE_LUT_B090 16'hB088
`define CUBE_LUT_B091 16'hB089
`define CUBE_LUT_B092 16'hB08A
`define CUBE_LUT_B093 16'hB08B
`define CUBE_LUT_B094 16'hB08C
`define CUBE_LUT_B095 16'hB08D
`define CUBE_LUT_B096 16'hB08E
`define CUBE_LUT_B097 16'hB08F
`define CUBE_LUT_B098 16'hB090
`define CUBE_LUT_B099 16'hB091
`define CUBE_LUT_B09A 16'hB092
`define CUBE_LUT_B09B 16'hB093
`define CUBE_LUT_B09C 16'hB094
`define CUBE_LUT_B09D 16'hB095
`define CUBE_LUT_B09E 16'hB096
`define CUBE_LUT_B09F 16'hB097
`define CUBE_LUT_B0A0 16'hB098
`define CUBE_LUT_B0A1 16'hB099
`define CUBE_LUT_B0A2 16'hB09A
`define CUBE_LUT_B0A3 16'hB09B
`define CUBE_LUT_B0A4 16'hB09C
`define CUBE_LUT_B0A5 16'hB09D
`define CUBE_LUT_B0A6 16'hB09E
`define CUBE_LUT_B0A7 16'hB09F
`define CUBE_LUT_B0A8 16'hB0A0
`define CUBE_LUT_B0A9 16'hB0A1
`define CUBE_LUT_B0AA 16'hB0A2
`define CUBE_LUT_B0AB 16'hB0A3
`define CUBE_LUT_B0AC 16'hB0A4
`define CUBE_LUT_B0AD 16'hB0A5
`define CUBE_LUT_B0AE 16'hB0A6
`define CUBE_LUT_B0AF 16'hB0A7
`define CUBE_LUT_B0B0 16'hB0A7
`define CUBE_LUT_B0B1 16'hB0A8
`define CUBE_LUT_B0B2 16'hB0A9
`define CUBE_LUT_B0B3 16'hB0AA
`define CUBE_LUT_B0B4 16'hB0AB
`define CUBE_LUT_B0B5 16'hB0AC
`define CUBE_LUT_B0B6 16'hB0AD
`define CUBE_LUT_B0B7 16'hB0AE
`define CUBE_LUT_B0B8 16'hB0AF
`define CUBE_LUT_B0B9 16'hB0B0
`define CUBE_LUT_B0BA 16'hB0B1
`define CUBE_LUT_B0BB 16'hB0B2
`define CUBE_LUT_B0BC 16'hB0B3
`define CUBE_LUT_B0BD 16'hB0B4
`define CUBE_LUT_B0BE 16'hB0B5
`define CUBE_LUT_B0BF 16'hB0B6
`define CUBE_LUT_B0C0 16'hB0B7
`define CUBE_LUT_B0C1 16'hB0B8
`define CUBE_LUT_B0C2 16'hB0B9
`define CUBE_LUT_B0C3 16'hB0BA
`define CUBE_LUT_B0C4 16'hB0BB
`define CUBE_LUT_B0C5 16'hB0BC
`define CUBE_LUT_B0C6 16'hB0BD
`define CUBE_LUT_B0C7 16'hB0BE
`define CUBE_LUT_B0C8 16'hB0BF
`define CUBE_LUT_B0C9 16'hB0C0
`define CUBE_LUT_B0CA 16'hB0C1
`define CUBE_LUT_B0CB 16'hB0C2
`define CUBE_LUT_B0CC 16'hB0C3
`define CUBE_LUT_B0CD 16'hB0C4
`define CUBE_LUT_B0CE 16'hB0C5
`define CUBE_LUT_B0CF 16'hB0C6
`define CUBE_LUT_B0D0 16'hB0C7
`define CUBE_LUT_B0D1 16'hB0C8
`define CUBE_LUT_B0D2 16'hB0C9
`define CUBE_LUT_B0D3 16'hB0CA
`define CUBE_LUT_B0D4 16'hB0CB
`define CUBE_LUT_B0D5 16'hB0CC
`define CUBE_LUT_B0D6 16'hB0CD
`define CUBE_LUT_B0D7 16'hB0CE
`define CUBE_LUT_B0D8 16'hB0CF
`define CUBE_LUT_B0D9 16'hB0D0
`define CUBE_LUT_B0DA 16'hB0D1
`define CUBE_LUT_B0DB 16'hB0D2
`define CUBE_LUT_B0DC 16'hB0D3
`define CUBE_LUT_B0DD 16'hB0D4
`define CUBE_LUT_B0DE 16'hB0D4
`define CUBE_LUT_B0DF 16'hB0D5
`define CUBE_LUT_B0E0 16'hB0D6
`define CUBE_LUT_B0E1 16'hB0D7
`define CUBE_LUT_B0E2 16'hB0D8
`define CUBE_LUT_B0E3 16'hB0D9
`define CUBE_LUT_B0E4 16'hB0DA
`define CUBE_LUT_B0E5 16'hB0DB
`define CUBE_LUT_B0E6 16'hB0DC
`define CUBE_LUT_B0E7 16'hB0DD
`define CUBE_LUT_B0E8 16'hB0DE
`define CUBE_LUT_B0E9 16'hB0DF
`define CUBE_LUT_B0EA 16'hB0E0
`define CUBE_LUT_B0EB 16'hB0E1
`define CUBE_LUT_B0EC 16'hB0E2
`define CUBE_LUT_B0ED 16'hB0E3
`define CUBE_LUT_B0EE 16'hB0E4
`define CUBE_LUT_B0EF 16'hB0E5
`define CUBE_LUT_B0F0 16'hB0E6
`define CUBE_LUT_B0F1 16'hB0E7
`define CUBE_LUT_B0F2 16'hB0E8
`define CUBE_LUT_B0F3 16'hB0E9
`define CUBE_LUT_B0F4 16'hB0EA
`define CUBE_LUT_B0F5 16'hB0EB
`define CUBE_LUT_B0F6 16'hB0EC
`define CUBE_LUT_B0F7 16'hB0ED
`define CUBE_LUT_B0F8 16'hB0EE
`define CUBE_LUT_B0F9 16'hB0EF
`define CUBE_LUT_B0FA 16'hB0F0
`define CUBE_LUT_B0FB 16'hB0F1
`define CUBE_LUT_B0FC 16'hB0F2
`define CUBE_LUT_B0FD 16'hB0F3
`define CUBE_LUT_B0FE 16'hB0F4
`define CUBE_LUT_B0FF 16'hB0F5
`define CUBE_LUT_B100 16'hB0F6
`define CUBE_LUT_B101 16'hB0F7
`define CUBE_LUT_B102 16'hB0F8
`define CUBE_LUT_B103 16'hB0F9
`define CUBE_LUT_B104 16'hB0FA
`define CUBE_LUT_B105 16'hB0FB
`define CUBE_LUT_B106 16'hB0FC
`define CUBE_LUT_B107 16'hB0FD
`define CUBE_LUT_B108 16'hB0FD
`define CUBE_LUT_B109 16'hB0FE
`define CUBE_LUT_B10A 16'hB0FF
`define CUBE_LUT_B10B 16'hB100
`define CUBE_LUT_B10C 16'hB101
`define CUBE_LUT_B10D 16'hB102
`define CUBE_LUT_B10E 16'hB103
`define CUBE_LUT_B10F 16'hB104
`define CUBE_LUT_B110 16'hB105
`define CUBE_LUT_B111 16'hB106
`define CUBE_LUT_B112 16'hB107
`define CUBE_LUT_B113 16'hB108
`define CUBE_LUT_B114 16'hB109
`define CUBE_LUT_B115 16'hB10A
`define CUBE_LUT_B116 16'hB10B
`define CUBE_LUT_B117 16'hB10C
`define CUBE_LUT_B118 16'hB10D
`define CUBE_LUT_B119 16'hB10E
`define CUBE_LUT_B11A 16'hB10F
`define CUBE_LUT_B11B 16'hB110
`define CUBE_LUT_B11C 16'hB111
`define CUBE_LUT_B11D 16'hB112
`define CUBE_LUT_B11E 16'hB113
`define CUBE_LUT_B11F 16'hB114
`define CUBE_LUT_B120 16'hB115
`define CUBE_LUT_B121 16'hB116
`define CUBE_LUT_B122 16'hB117
`define CUBE_LUT_B123 16'hB118
`define CUBE_LUT_B124 16'hB119
`define CUBE_LUT_B125 16'hB11A
`define CUBE_LUT_B126 16'hB11B
`define CUBE_LUT_B127 16'hB11C
`define CUBE_LUT_B128 16'hB11D
`define CUBE_LUT_B129 16'hB11E
`define CUBE_LUT_B12A 16'hB11F
`define CUBE_LUT_B12B 16'hB120
`define CUBE_LUT_B12C 16'hB121
`define CUBE_LUT_B12D 16'hB122
`define CUBE_LUT_B12E 16'hB123
`define CUBE_LUT_B12F 16'hB124
`define CUBE_LUT_B130 16'hB124
`define CUBE_LUT_B131 16'hB125
`define CUBE_LUT_B132 16'hB126
`define CUBE_LUT_B133 16'hB127
`define CUBE_LUT_B134 16'hB128
`define CUBE_LUT_B135 16'hB129
`define CUBE_LUT_B136 16'hB12A
`define CUBE_LUT_B137 16'hB12B
`define CUBE_LUT_B138 16'hB12C
`define CUBE_LUT_B139 16'hB12D
`define CUBE_LUT_B13A 16'hB12E
`define CUBE_LUT_B13B 16'hB12F
`define CUBE_LUT_B13C 16'hB130
`define CUBE_LUT_B13D 16'hB131
`define CUBE_LUT_B13E 16'hB132
`define CUBE_LUT_B13F 16'hB133
`define CUBE_LUT_B140 16'hB134
`define CUBE_LUT_B141 16'hB135
`define CUBE_LUT_B142 16'hB136
`define CUBE_LUT_B143 16'hB137
`define CUBE_LUT_B144 16'hB138
`define CUBE_LUT_B145 16'hB139
`define CUBE_LUT_B146 16'hB13A
`define CUBE_LUT_B147 16'hB13B
`define CUBE_LUT_B148 16'hB13C
`define CUBE_LUT_B149 16'hB13D
`define CUBE_LUT_B14A 16'hB13E
`define CUBE_LUT_B14B 16'hB13F
`define CUBE_LUT_B14C 16'hB140
`define CUBE_LUT_B14D 16'hB141
`define CUBE_LUT_B14E 16'hB142
`define CUBE_LUT_B14F 16'hB143
`define CUBE_LUT_B150 16'hB144
`define CUBE_LUT_B151 16'hB145
`define CUBE_LUT_B152 16'hB146
`define CUBE_LUT_B153 16'hB147
`define CUBE_LUT_B154 16'hB148
`define CUBE_LUT_B155 16'hB149
`define CUBE_LUT_B156 16'hB149
`define CUBE_LUT_B157 16'hB14A
`define CUBE_LUT_B158 16'hB14B
`define CUBE_LUT_B159 16'hB14C
`define CUBE_LUT_B15A 16'hB14D
`define CUBE_LUT_B15B 16'hB14E
`define CUBE_LUT_B15C 16'hB14F
`define CUBE_LUT_B15D 16'hB150
`define CUBE_LUT_B15E 16'hB151
`define CUBE_LUT_B15F 16'hB152
`define CUBE_LUT_B160 16'hB153
`define CUBE_LUT_B161 16'hB154
`define CUBE_LUT_B162 16'hB155
`define CUBE_LUT_B163 16'hB156
`define CUBE_LUT_B164 16'hB157
`define CUBE_LUT_B165 16'hB158
`define CUBE_LUT_B166 16'hB159
`define CUBE_LUT_B167 16'hB15A
`define CUBE_LUT_B168 16'hB15B
`define CUBE_LUT_B169 16'hB15C
`define CUBE_LUT_B16A 16'hB15D
`define CUBE_LUT_B16B 16'hB15E
`define CUBE_LUT_B16C 16'hB15F
`define CUBE_LUT_B16D 16'hB160
`define CUBE_LUT_B16E 16'hB161
`define CUBE_LUT_B16F 16'hB162
`define CUBE_LUT_B170 16'hB163
`define CUBE_LUT_B171 16'hB164
`define CUBE_LUT_B172 16'hB165
`define CUBE_LUT_B173 16'hB166
`define CUBE_LUT_B174 16'hB167
`define CUBE_LUT_B175 16'hB168
`define CUBE_LUT_B176 16'hB169
`define CUBE_LUT_B177 16'hB16A
`define CUBE_LUT_B178 16'hB16B
`define CUBE_LUT_B179 16'hB16B
`define CUBE_LUT_B17A 16'hB16C
`define CUBE_LUT_B17B 16'hB16D
`define CUBE_LUT_B17C 16'hB16E
`define CUBE_LUT_B17D 16'hB16F
`define CUBE_LUT_B17E 16'hB170
`define CUBE_LUT_B17F 16'hB171
`define CUBE_LUT_B180 16'hB172
`define CUBE_LUT_B181 16'hB173
`define CUBE_LUT_B182 16'hB174
`define CUBE_LUT_B183 16'hB175
`define CUBE_LUT_B184 16'hB176
`define CUBE_LUT_B185 16'hB177
`define CUBE_LUT_B186 16'hB178
`define CUBE_LUT_B187 16'hB179
`define CUBE_LUT_B188 16'hB17A
`define CUBE_LUT_B189 16'hB17B
`define CUBE_LUT_B18A 16'hB17C
`define CUBE_LUT_B18B 16'hB17D
`define CUBE_LUT_B18C 16'hB17E
`define CUBE_LUT_B18D 16'hB17F
`define CUBE_LUT_B18E 16'hB180
`define CUBE_LUT_B18F 16'hB181
`define CUBE_LUT_B190 16'hB182
`define CUBE_LUT_B191 16'hB183
`define CUBE_LUT_B192 16'hB184
`define CUBE_LUT_B193 16'hB185
`define CUBE_LUT_B194 16'hB186
`define CUBE_LUT_B195 16'hB187
`define CUBE_LUT_B196 16'hB188
`define CUBE_LUT_B197 16'hB189
`define CUBE_LUT_B198 16'hB18A
`define CUBE_LUT_B199 16'hB18B
`define CUBE_LUT_B19A 16'hB18C
`define CUBE_LUT_B19B 16'hB18D
`define CUBE_LUT_B19C 16'hB18D
`define CUBE_LUT_B19D 16'hB18E
`define CUBE_LUT_B19E 16'hB18F
`define CUBE_LUT_B19F 16'hB190
`define CUBE_LUT_B1A0 16'hB191
`define CUBE_LUT_B1A1 16'hB192
`define CUBE_LUT_B1A2 16'hB193
`define CUBE_LUT_B1A3 16'hB194
`define CUBE_LUT_B1A4 16'hB195
`define CUBE_LUT_B1A5 16'hB196
`define CUBE_LUT_B1A6 16'hB197
`define CUBE_LUT_B1A7 16'hB198
`define CUBE_LUT_B1A8 16'hB199
`define CUBE_LUT_B1A9 16'hB19A
`define CUBE_LUT_B1AA 16'hB19B
`define CUBE_LUT_B1AB 16'hB19C
`define CUBE_LUT_B1AC 16'hB19D
`define CUBE_LUT_B1AD 16'hB19E
`define CUBE_LUT_B1AE 16'hB19F
`define CUBE_LUT_B1AF 16'hB1A0
`define CUBE_LUT_B1B0 16'hB1A1
`define CUBE_LUT_B1B1 16'hB1A2
`define CUBE_LUT_B1B2 16'hB1A3
`define CUBE_LUT_B1B3 16'hB1A4
`define CUBE_LUT_B1B4 16'hB1A5
`define CUBE_LUT_B1B5 16'hB1A6
`define CUBE_LUT_B1B6 16'hB1A7
`define CUBE_LUT_B1B7 16'hB1A8
`define CUBE_LUT_B1B8 16'hB1A9
`define CUBE_LUT_B1B9 16'hB1AA
`define CUBE_LUT_B1BA 16'hB1AB
`define CUBE_LUT_B1BB 16'hB1AC
`define CUBE_LUT_B1BC 16'hB1AC
`define CUBE_LUT_B1BD 16'hB1AD
`define CUBE_LUT_B1BE 16'hB1AE
`define CUBE_LUT_B1BF 16'hB1AF
`define CUBE_LUT_B1C0 16'hB1B0
`define CUBE_LUT_B1C1 16'hB1B1
`define CUBE_LUT_B1C2 16'hB1B2
`define CUBE_LUT_B1C3 16'hB1B3
`define CUBE_LUT_B1C4 16'hB1B4
`define CUBE_LUT_B1C5 16'hB1B5
`define CUBE_LUT_B1C6 16'hB1B6
`define CUBE_LUT_B1C7 16'hB1B7
`define CUBE_LUT_B1C8 16'hB1B8
`define CUBE_LUT_B1C9 16'hB1B9
`define CUBE_LUT_B1CA 16'hB1BA
`define CUBE_LUT_B1CB 16'hB1BB
`define CUBE_LUT_B1CC 16'hB1BC
`define CUBE_LUT_B1CD 16'hB1BD
`define CUBE_LUT_B1CE 16'hB1BE
`define CUBE_LUT_B1CF 16'hB1BF
`define CUBE_LUT_B1D0 16'hB1C0
`define CUBE_LUT_B1D1 16'hB1C1
`define CUBE_LUT_B1D2 16'hB1C2
`define CUBE_LUT_B1D3 16'hB1C3
`define CUBE_LUT_B1D4 16'hB1C4
`define CUBE_LUT_B1D5 16'hB1C5
`define CUBE_LUT_B1D6 16'hB1C6
`define CUBE_LUT_B1D7 16'hB1C7
`define CUBE_LUT_B1D8 16'hB1C8
`define CUBE_LUT_B1D9 16'hB1C9
`define CUBE_LUT_B1DA 16'hB1CA
`define CUBE_LUT_B1DB 16'hB1CA
`define CUBE_LUT_B1DC 16'hB1CB
`define CUBE_LUT_B1DD 16'hB1CC
`define CUBE_LUT_B1DE 16'hB1CD
`define CUBE_LUT_B1DF 16'hB1CE
`define CUBE_LUT_B1E0 16'hB1CF
`define CUBE_LUT_B1E1 16'hB1D0
`define CUBE_LUT_B1E2 16'hB1D1
`define CUBE_LUT_B1E3 16'hB1D2
`define CUBE_LUT_B1E4 16'hB1D3
`define CUBE_LUT_B1E5 16'hB1D4
`define CUBE_LUT_B1E6 16'hB1D5
`define CUBE_LUT_B1E7 16'hB1D6
`define CUBE_LUT_B1E8 16'hB1D7
`define CUBE_LUT_B1E9 16'hB1D8
`define CUBE_LUT_B1EA 16'hB1D9
`define CUBE_LUT_B1EB 16'hB1DA
`define CUBE_LUT_B1EC 16'hB1DB
`define CUBE_LUT_B1ED 16'hB1DC
`define CUBE_LUT_B1EE 16'hB1DD
`define CUBE_LUT_B1EF 16'hB1DE
`define CUBE_LUT_B1F0 16'hB1DF
`define CUBE_LUT_B1F1 16'hB1E0
`define CUBE_LUT_B1F2 16'hB1E1
`define CUBE_LUT_B1F3 16'hB1E2
`define CUBE_LUT_B1F4 16'hB1E3
`define CUBE_LUT_B1F5 16'hB1E4
`define CUBE_LUT_B1F6 16'hB1E5
`define CUBE_LUT_B1F7 16'hB1E6
`define CUBE_LUT_B1F8 16'hB1E7
`define CUBE_LUT_B1F9 16'hB1E7
`define CUBE_LUT_B1FA 16'hB1E8
`define CUBE_LUT_B1FB 16'hB1E9
`define CUBE_LUT_B1FC 16'hB1EA
`define CUBE_LUT_B1FD 16'hB1EB
`define CUBE_LUT_B1FE 16'hB1EC
`define CUBE_LUT_B1FF 16'hB1ED
`define CUBE_LUT_B200 16'hB1EE
`define CUBE_LUT_B201 16'hB1EF
`define CUBE_LUT_B202 16'hB1F0
`define CUBE_LUT_B203 16'hB1F1
`define CUBE_LUT_B204 16'hB1F2
`define CUBE_LUT_B205 16'hB1F3
`define CUBE_LUT_B206 16'hB1F4
`define CUBE_LUT_B207 16'hB1F5
`define CUBE_LUT_B208 16'hB1F6
`define CUBE_LUT_B209 16'hB1F7
`define CUBE_LUT_B20A 16'hB1F8
`define CUBE_LUT_B20B 16'hB1F9
`define CUBE_LUT_B20C 16'hB1FA
`define CUBE_LUT_B20D 16'hB1FB
`define CUBE_LUT_B20E 16'hB1FC
`define CUBE_LUT_B20F 16'hB1FD
`define CUBE_LUT_B210 16'hB1FE
`define CUBE_LUT_B211 16'hB1FF
`define CUBE_LUT_B212 16'hB200
`define CUBE_LUT_B213 16'hB201
`define CUBE_LUT_B214 16'hB202
`define CUBE_LUT_B215 16'hB203
`define CUBE_LUT_B216 16'hB203
`define CUBE_LUT_B217 16'hB204
`define CUBE_LUT_B218 16'hB205
`define CUBE_LUT_B219 16'hB206
`define CUBE_LUT_B21A 16'hB207
`define CUBE_LUT_B21B 16'hB208
`define CUBE_LUT_B21C 16'hB209
`define CUBE_LUT_B21D 16'hB20A
`define CUBE_LUT_B21E 16'hB20B
`define CUBE_LUT_B21F 16'hB20C
`define CUBE_LUT_B220 16'hB20D
`define CUBE_LUT_B221 16'hB20E
`define CUBE_LUT_B222 16'hB20F
`define CUBE_LUT_B223 16'hB210
`define CUBE_LUT_B224 16'hB211
`define CUBE_LUT_B225 16'hB212
`define CUBE_LUT_B226 16'hB213
`define CUBE_LUT_B227 16'hB214
`define CUBE_LUT_B228 16'hB215
`define CUBE_LUT_B229 16'hB216
`define CUBE_LUT_B22A 16'hB217
`define CUBE_LUT_B22B 16'hB218
`define CUBE_LUT_B22C 16'hB219
`define CUBE_LUT_B22D 16'hB21A
`define CUBE_LUT_B22E 16'hB21B
`define CUBE_LUT_B22F 16'hB21C
`define CUBE_LUT_B230 16'hB21D
`define CUBE_LUT_B231 16'hB21E
`define CUBE_LUT_B232 16'hB21E
`define CUBE_LUT_B233 16'hB21F
`define CUBE_LUT_B234 16'hB220
`define CUBE_LUT_B235 16'hB221
`define CUBE_LUT_B236 16'hB222
`define CUBE_LUT_B237 16'hB223
`define CUBE_LUT_B238 16'hB224
`define CUBE_LUT_B239 16'hB225
`define CUBE_LUT_B23A 16'hB226
`define CUBE_LUT_B23B 16'hB227
`define CUBE_LUT_B23C 16'hB228
`define CUBE_LUT_B23D 16'hB229
`define CUBE_LUT_B23E 16'hB22A
`define CUBE_LUT_B23F 16'hB22B
`define CUBE_LUT_B240 16'hB22C
`define CUBE_LUT_B241 16'hB22D
`define CUBE_LUT_B242 16'hB22E
`define CUBE_LUT_B243 16'hB22F
`define CUBE_LUT_B244 16'hB230
`define CUBE_LUT_B245 16'hB231
`define CUBE_LUT_B246 16'hB232
`define CUBE_LUT_B247 16'hB233
`define CUBE_LUT_B248 16'hB234
`define CUBE_LUT_B249 16'hB235
`define CUBE_LUT_B24A 16'hB236
`define CUBE_LUT_B24B 16'hB237
`define CUBE_LUT_B24C 16'hB238
`define CUBE_LUT_B24D 16'hB238
`define CUBE_LUT_B24E 16'hB239
`define CUBE_LUT_B24F 16'hB23A
`define CUBE_LUT_B250 16'hB23B
`define CUBE_LUT_B251 16'hB23C
`define CUBE_LUT_B252 16'hB23D
`define CUBE_LUT_B253 16'hB23E
`define CUBE_LUT_B254 16'hB23F
`define CUBE_LUT_B255 16'hB240
`define CUBE_LUT_B256 16'hB241
`define CUBE_LUT_B257 16'hB242
`define CUBE_LUT_B258 16'hB243
`define CUBE_LUT_B259 16'hB244
`define CUBE_LUT_B25A 16'hB245
`define CUBE_LUT_B25B 16'hB246
`define CUBE_LUT_B25C 16'hB247
`define CUBE_LUT_B25D 16'hB248
`define CUBE_LUT_B25E 16'hB249
`define CUBE_LUT_B25F 16'hB24A
`define CUBE_LUT_B260 16'hB24B
`define CUBE_LUT_B261 16'hB24C
`define CUBE_LUT_B262 16'hB24D
`define CUBE_LUT_B263 16'hB24E
`define CUBE_LUT_B264 16'hB24F
`define CUBE_LUT_B265 16'hB250
`define CUBE_LUT_B266 16'hB251
`define CUBE_LUT_B267 16'hB251
`define CUBE_LUT_B268 16'hB252
`define CUBE_LUT_B269 16'hB253
`define CUBE_LUT_B26A 16'hB254
`define CUBE_LUT_B26B 16'hB255
`define CUBE_LUT_B26C 16'hB256
`define CUBE_LUT_B26D 16'hB257
`define CUBE_LUT_B26E 16'hB258
`define CUBE_LUT_B26F 16'hB259
`define CUBE_LUT_B270 16'hB25A
`define CUBE_LUT_B271 16'hB25B
`define CUBE_LUT_B272 16'hB25C
`define CUBE_LUT_B273 16'hB25D
`define CUBE_LUT_B274 16'hB25E
`define CUBE_LUT_B275 16'hB25F
`define CUBE_LUT_B276 16'hB260
`define CUBE_LUT_B277 16'hB261
`define CUBE_LUT_B278 16'hB262
`define CUBE_LUT_B279 16'hB263
`define CUBE_LUT_B27A 16'hB264
`define CUBE_LUT_B27B 16'hB265
`define CUBE_LUT_B27C 16'hB266
`define CUBE_LUT_B27D 16'hB267
`define CUBE_LUT_B27E 16'hB268
`define CUBE_LUT_B27F 16'hB269
`define CUBE_LUT_B280 16'hB269
`define CUBE_LUT_B281 16'hB26A
`define CUBE_LUT_B282 16'hB26B
`define CUBE_LUT_B283 16'hB26C
`define CUBE_LUT_B284 16'hB26D
`define CUBE_LUT_B285 16'hB26E
`define CUBE_LUT_B286 16'hB26F
`define CUBE_LUT_B287 16'hB270
`define CUBE_LUT_B288 16'hB271
`define CUBE_LUT_B289 16'hB272
`define CUBE_LUT_B28A 16'hB273
`define CUBE_LUT_B28B 16'hB274
`define CUBE_LUT_B28C 16'hB275
`define CUBE_LUT_B28D 16'hB276
`define CUBE_LUT_B28E 16'hB277
`define CUBE_LUT_B28F 16'hB278
`define CUBE_LUT_B290 16'hB279
`define CUBE_LUT_B291 16'hB27A
`define CUBE_LUT_B292 16'hB27B
`define CUBE_LUT_B293 16'hB27C
`define CUBE_LUT_B294 16'hB27D
`define CUBE_LUT_B295 16'hB27E
`define CUBE_LUT_B296 16'hB27F
`define CUBE_LUT_B297 16'hB280
`define CUBE_LUT_B298 16'hB281
`define CUBE_LUT_B299 16'hB281
`define CUBE_LUT_B29A 16'hB282
`define CUBE_LUT_B29B 16'hB283
`define CUBE_LUT_B29C 16'hB284
`define CUBE_LUT_B29D 16'hB285
`define CUBE_LUT_B29E 16'hB286
`define CUBE_LUT_B29F 16'hB287
`define CUBE_LUT_B2A0 16'hB288
`define CUBE_LUT_B2A1 16'hB289
`define CUBE_LUT_B2A2 16'hB28A
`define CUBE_LUT_B2A3 16'hB28B
`define CUBE_LUT_B2A4 16'hB28C
`define CUBE_LUT_B2A5 16'hB28D
`define CUBE_LUT_B2A6 16'hB28E
`define CUBE_LUT_B2A7 16'hB28F
`define CUBE_LUT_B2A8 16'hB290
`define CUBE_LUT_B2A9 16'hB291
`define CUBE_LUT_B2AA 16'hB292
`define CUBE_LUT_B2AB 16'hB293
`define CUBE_LUT_B2AC 16'hB294
`define CUBE_LUT_B2AD 16'hB295
`define CUBE_LUT_B2AE 16'hB296
`define CUBE_LUT_B2AF 16'hB297
`define CUBE_LUT_B2B0 16'hB298
`define CUBE_LUT_B2B1 16'hB298
`define CUBE_LUT_B2B2 16'hB299
`define CUBE_LUT_B2B3 16'hB29A
`define CUBE_LUT_B2B4 16'hB29B
`define CUBE_LUT_B2B5 16'hB29C
`define CUBE_LUT_B2B6 16'hB29D
`define CUBE_LUT_B2B7 16'hB29E
`define CUBE_LUT_B2B8 16'hB29F
`define CUBE_LUT_B2B9 16'hB2A0
`define CUBE_LUT_B2BA 16'hB2A1
`define CUBE_LUT_B2BB 16'hB2A2
`define CUBE_LUT_B2BC 16'hB2A3
`define CUBE_LUT_B2BD 16'hB2A4
`define CUBE_LUT_B2BE 16'hB2A5
`define CUBE_LUT_B2BF 16'hB2A6
`define CUBE_LUT_B2C0 16'hB2A7
`define CUBE_LUT_B2C1 16'hB2A8
`define CUBE_LUT_B2C2 16'hB2A9
`define CUBE_LUT_B2C3 16'hB2AA
`define CUBE_LUT_B2C4 16'hB2AB
`define CUBE_LUT_B2C5 16'hB2AC
`define CUBE_LUT_B2C6 16'hB2AD
`define CUBE_LUT_B2C7 16'hB2AE
`define CUBE_LUT_B2C8 16'hB2AE
`define CUBE_LUT_B2C9 16'hB2AF
`define CUBE_LUT_B2CA 16'hB2B0
`define CUBE_LUT_B2CB 16'hB2B1
`define CUBE_LUT_B2CC 16'hB2B2
`define CUBE_LUT_B2CD 16'hB2B3
`define CUBE_LUT_B2CE 16'hB2B4
`define CUBE_LUT_B2CF 16'hB2B5
`define CUBE_LUT_B2D0 16'hB2B6
`define CUBE_LUT_B2D1 16'hB2B7
`define CUBE_LUT_B2D2 16'hB2B8
`define CUBE_LUT_B2D3 16'hB2B9
`define CUBE_LUT_B2D4 16'hB2BA
`define CUBE_LUT_B2D5 16'hB2BB
`define CUBE_LUT_B2D6 16'hB2BC
`define CUBE_LUT_B2D7 16'hB2BD
`define CUBE_LUT_B2D8 16'hB2BE
`define CUBE_LUT_B2D9 16'hB2BF
`define CUBE_LUT_B2DA 16'hB2C0
`define CUBE_LUT_B2DB 16'hB2C1
`define CUBE_LUT_B2DC 16'hB2C2
`define CUBE_LUT_B2DD 16'hB2C3
`define CUBE_LUT_B2DE 16'hB2C4
`define CUBE_LUT_B2DF 16'hB2C4
`define CUBE_LUT_B2E0 16'hB2C5
`define CUBE_LUT_B2E1 16'hB2C6
`define CUBE_LUT_B2E2 16'hB2C7
`define CUBE_LUT_B2E3 16'hB2C8
`define CUBE_LUT_B2E4 16'hB2C9
`define CUBE_LUT_B2E5 16'hB2CA
`define CUBE_LUT_B2E6 16'hB2CB
`define CUBE_LUT_B2E7 16'hB2CC
`define CUBE_LUT_B2E8 16'hB2CD
`define CUBE_LUT_B2E9 16'hB2CE
`define CUBE_LUT_B2EA 16'hB2CF
`define CUBE_LUT_B2EB 16'hB2D0
`define CUBE_LUT_B2EC 16'hB2D1
`define CUBE_LUT_B2ED 16'hB2D2
`define CUBE_LUT_B2EE 16'hB2D3
`define CUBE_LUT_B2EF 16'hB2D4
`define CUBE_LUT_B2F0 16'hB2D5
`define CUBE_LUT_B2F1 16'hB2D6
`define CUBE_LUT_B2F2 16'hB2D7
`define CUBE_LUT_B2F3 16'hB2D8
`define CUBE_LUT_B2F4 16'hB2D9
`define CUBE_LUT_B2F5 16'hB2D9
`define CUBE_LUT_B2F6 16'hB2DA
`define CUBE_LUT_B2F7 16'hB2DB
`define CUBE_LUT_B2F8 16'hB2DC
`define CUBE_LUT_B2F9 16'hB2DD
`define CUBE_LUT_B2FA 16'hB2DE
`define CUBE_LUT_B2FB 16'hB2DF
`define CUBE_LUT_B2FC 16'hB2E0
`define CUBE_LUT_B2FD 16'hB2E1
`define CUBE_LUT_B2FE 16'hB2E2
`define CUBE_LUT_B2FF 16'hB2E3
`define CUBE_LUT_B300 16'hB2E4
`define CUBE_LUT_B301 16'hB2E5
`define CUBE_LUT_B302 16'hB2E6
`define CUBE_LUT_B303 16'hB2E7
`define CUBE_LUT_B304 16'hB2E8
`define CUBE_LUT_B305 16'hB2E9
`define CUBE_LUT_B306 16'hB2EA
`define CUBE_LUT_B307 16'hB2EB
`define CUBE_LUT_B308 16'hB2EC
`define CUBE_LUT_B309 16'hB2ED
`define CUBE_LUT_B30A 16'hB2ED
`define CUBE_LUT_B30B 16'hB2EE
`define CUBE_LUT_B30C 16'hB2EF
`define CUBE_LUT_B30D 16'hB2F0
`define CUBE_LUT_B30E 16'hB2F1
`define CUBE_LUT_B30F 16'hB2F2
`define CUBE_LUT_B310 16'hB2F3
`define CUBE_LUT_B311 16'hB2F4
`define CUBE_LUT_B312 16'hB2F5
`define CUBE_LUT_B313 16'hB2F6
`define CUBE_LUT_B314 16'hB2F7
`define CUBE_LUT_B315 16'hB2F8
`define CUBE_LUT_B316 16'hB2F9
`define CUBE_LUT_B317 16'hB2FA
`define CUBE_LUT_B318 16'hB2FB
`define CUBE_LUT_B319 16'hB2FC
`define CUBE_LUT_B31A 16'hB2FD
`define CUBE_LUT_B31B 16'hB2FE
`define CUBE_LUT_B31C 16'hB2FF
`define CUBE_LUT_B31D 16'hB300
`define CUBE_LUT_B31E 16'hB301
`define CUBE_LUT_B31F 16'hB301
`define CUBE_LUT_B320 16'hB302
`define CUBE_LUT_B321 16'hB303
`define CUBE_LUT_B322 16'hB304
`define CUBE_LUT_B323 16'hB305
`define CUBE_LUT_B324 16'hB306
`define CUBE_LUT_B325 16'hB307
`define CUBE_LUT_B326 16'hB308
`define CUBE_LUT_B327 16'hB309
`define CUBE_LUT_B328 16'hB30A
`define CUBE_LUT_B329 16'hB30B
`define CUBE_LUT_B32A 16'hB30C
`define CUBE_LUT_B32B 16'hB30D
`define CUBE_LUT_B32C 16'hB30E
`define CUBE_LUT_B32D 16'hB30F
`define CUBE_LUT_B32E 16'hB310
`define CUBE_LUT_B32F 16'hB311
`define CUBE_LUT_B330 16'hB312
`define CUBE_LUT_B331 16'hB313
`define CUBE_LUT_B332 16'hB314
`define CUBE_LUT_B333 16'hB315
`define CUBE_LUT_B334 16'hB315
`define CUBE_LUT_B335 16'hB316
`define CUBE_LUT_B336 16'hB317
`define CUBE_LUT_B337 16'hB318
`define CUBE_LUT_B338 16'hB319
`define CUBE_LUT_B339 16'hB31A
`define CUBE_LUT_B33A 16'hB31B
`define CUBE_LUT_B33B 16'hB31C
`define CUBE_LUT_B33C 16'hB31D
`define CUBE_LUT_B33D 16'hB31E
`define CUBE_LUT_B33E 16'hB31F
`define CUBE_LUT_B33F 16'hB320
`define CUBE_LUT_B340 16'hB321
`define CUBE_LUT_B341 16'hB322
`define CUBE_LUT_B342 16'hB323
`define CUBE_LUT_B343 16'hB324
`define CUBE_LUT_B344 16'hB325
`define CUBE_LUT_B345 16'hB326
`define CUBE_LUT_B346 16'hB327
`define CUBE_LUT_B347 16'hB328
`define CUBE_LUT_B348 16'hB328
`define CUBE_LUT_B349 16'hB329
`define CUBE_LUT_B34A 16'hB32A
`define CUBE_LUT_B34B 16'hB32B
`define CUBE_LUT_B34C 16'hB32C
`define CUBE_LUT_B34D 16'hB32D
`define CUBE_LUT_B34E 16'hB32E
`define CUBE_LUT_B34F 16'hB32F
`define CUBE_LUT_B350 16'hB330
`define CUBE_LUT_B351 16'hB331
`define CUBE_LUT_B352 16'hB332
`define CUBE_LUT_B353 16'hB333
`define CUBE_LUT_B354 16'hB334
`define CUBE_LUT_B355 16'hB335
`define CUBE_LUT_B356 16'hB336
`define CUBE_LUT_B357 16'hB337
`define CUBE_LUT_B358 16'hB338
`define CUBE_LUT_B359 16'hB339
`define CUBE_LUT_B35A 16'hB33A
`define CUBE_LUT_B35B 16'hB33B
`define CUBE_LUT_B35C 16'hB33B
`define CUBE_LUT_B35D 16'hB33C
`define CUBE_LUT_B35E 16'hB33D
`define CUBE_LUT_B35F 16'hB33E
`define CUBE_LUT_B360 16'hB33F
`define CUBE_LUT_B361 16'hB340
`define CUBE_LUT_B362 16'hB341
`define CUBE_LUT_B363 16'hB342
`define CUBE_LUT_B364 16'hB343
`define CUBE_LUT_B365 16'hB344
`define CUBE_LUT_B366 16'hB345
`define CUBE_LUT_B367 16'hB346
`define CUBE_LUT_B368 16'hB347
`define CUBE_LUT_B369 16'hB348
`define CUBE_LUT_B36A 16'hB349
`define CUBE_LUT_B36B 16'hB34A
`define CUBE_LUT_B36C 16'hB34B
`define CUBE_LUT_B36D 16'hB34C
`define CUBE_LUT_B36E 16'hB34D
`define CUBE_LUT_B36F 16'hB34D
`define CUBE_LUT_B370 16'hB34E
`define CUBE_LUT_B371 16'hB34F
`define CUBE_LUT_B372 16'hB350
`define CUBE_LUT_B373 16'hB351
`define CUBE_LUT_B374 16'hB352
`define CUBE_LUT_B375 16'hB353
`define CUBE_LUT_B376 16'hB354
`define CUBE_LUT_B377 16'hB355
`define CUBE_LUT_B378 16'hB356
`define CUBE_LUT_B379 16'hB357
`define CUBE_LUT_B37A 16'hB358
`define CUBE_LUT_B37B 16'hB359
`define CUBE_LUT_B37C 16'hB35A
`define CUBE_LUT_B37D 16'hB35B
`define CUBE_LUT_B37E 16'hB35C
`define CUBE_LUT_B37F 16'hB35D
`define CUBE_LUT_B380 16'hB35E
`define CUBE_LUT_B381 16'hB35F
`define CUBE_LUT_B382 16'hB35F
`define CUBE_LUT_B383 16'hB360
`define CUBE_LUT_B384 16'hB361
`define CUBE_LUT_B385 16'hB362
`define CUBE_LUT_B386 16'hB363
`define CUBE_LUT_B387 16'hB364
`define CUBE_LUT_B388 16'hB365
`define CUBE_LUT_B389 16'hB366
`define CUBE_LUT_B38A 16'hB367
`define CUBE_LUT_B38B 16'hB368
`define CUBE_LUT_B38C 16'hB369
`define CUBE_LUT_B38D 16'hB36A
`define CUBE_LUT_B38E 16'hB36B
`define CUBE_LUT_B38F 16'hB36C
`define CUBE_LUT_B390 16'hB36D
`define CUBE_LUT_B391 16'hB36E
`define CUBE_LUT_B392 16'hB36F
`define CUBE_LUT_B393 16'hB370
`define CUBE_LUT_B394 16'hB371
`define CUBE_LUT_B395 16'hB371
`define CUBE_LUT_B396 16'hB372
`define CUBE_LUT_B397 16'hB373
`define CUBE_LUT_B398 16'hB374
`define CUBE_LUT_B399 16'hB375
`define CUBE_LUT_B39A 16'hB376
`define CUBE_LUT_B39B 16'hB377
`define CUBE_LUT_B39C 16'hB378
`define CUBE_LUT_B39D 16'hB379
`define CUBE_LUT_B39E 16'hB37A
`define CUBE_LUT_B39F 16'hB37B
`define CUBE_LUT_B3A0 16'hB37C
`define CUBE_LUT_B3A1 16'hB37D
`define CUBE_LUT_B3A2 16'hB37E
`define CUBE_LUT_B3A3 16'hB37F
`define CUBE_LUT_B3A4 16'hB380
`define CUBE_LUT_B3A5 16'hB381
`define CUBE_LUT_B3A6 16'hB382
`define CUBE_LUT_B3A7 16'hB382
`define CUBE_LUT_B3A8 16'hB383
`define CUBE_LUT_B3A9 16'hB384
`define CUBE_LUT_B3AA 16'hB385
`define CUBE_LUT_B3AB 16'hB386
`define CUBE_LUT_B3AC 16'hB387
`define CUBE_LUT_B3AD 16'hB388
`define CUBE_LUT_B3AE 16'hB389
`define CUBE_LUT_B3AF 16'hB38A
`define CUBE_LUT_B3B0 16'hB38B
`define CUBE_LUT_B3B1 16'hB38C
`define CUBE_LUT_B3B2 16'hB38D
`define CUBE_LUT_B3B3 16'hB38E
`define CUBE_LUT_B3B4 16'hB38F
`define CUBE_LUT_B3B5 16'hB390
`define CUBE_LUT_B3B6 16'hB391
`define CUBE_LUT_B3B7 16'hB392
`define CUBE_LUT_B3B8 16'hB393
`define CUBE_LUT_B3B9 16'hB393
`define CUBE_LUT_B3BA 16'hB394
`define CUBE_LUT_B3BB 16'hB395
`define CUBE_LUT_B3BC 16'hB396
`define CUBE_LUT_B3BD 16'hB397
`define CUBE_LUT_B3BE 16'hB398
`define CUBE_LUT_B3BF 16'hB399
`define CUBE_LUT_B3C0 16'hB39A
`define CUBE_LUT_B3C1 16'hB39B
`define CUBE_LUT_B3C2 16'hB39C
`define CUBE_LUT_B3C3 16'hB39D
`define CUBE_LUT_B3C4 16'hB39E
`define CUBE_LUT_B3C5 16'hB39F
`define CUBE_LUT_B3C6 16'hB3A0
`define CUBE_LUT_B3C7 16'hB3A1
`define CUBE_LUT_B3C8 16'hB3A2
`define CUBE_LUT_B3C9 16'hB3A3
`define CUBE_LUT_B3CA 16'hB3A4
`define CUBE_LUT_B3CB 16'hB3A4
`define CUBE_LUT_B3CC 16'hB3A5
`define CUBE_LUT_B3CD 16'hB3A6
`define CUBE_LUT_B3CE 16'hB3A7
`define CUBE_LUT_B3CF 16'hB3A8
`define CUBE_LUT_B3D0 16'hB3A9
`define CUBE_LUT_B3D1 16'hB3AA
`define CUBE_LUT_B3D2 16'hB3AB
`define CUBE_LUT_B3D3 16'hB3AC
`define CUBE_LUT_B3D4 16'hB3AD
`define CUBE_LUT_B3D5 16'hB3AE
`define CUBE_LUT_B3D6 16'hB3AF
`define CUBE_LUT_B3D7 16'hB3B0
`define CUBE_LUT_B3D8 16'hB3B1
`define CUBE_LUT_B3D9 16'hB3B2
`define CUBE_LUT_B3DA 16'hB3B3
`define CUBE_LUT_B3DB 16'hB3B4
`define CUBE_LUT_B3DC 16'hB3B4
`define CUBE_LUT_B3DD 16'hB3B5
`define CUBE_LUT_B3DE 16'hB3B6
`define CUBE_LUT_B3DF 16'hB3B7
`define CUBE_LUT_B3E0 16'hB3B8
`define CUBE_LUT_B3E1 16'hB3B9
`define CUBE_LUT_B3E2 16'hB3BA
`define CUBE_LUT_B3E3 16'hB3BB
`define CUBE_LUT_B3E4 16'hB3BC
`define CUBE_LUT_B3E5 16'hB3BD
`define CUBE_LUT_B3E6 16'hB3BE
`define CUBE_LUT_B3E7 16'hB3BF
`define CUBE_LUT_B3E8 16'hB3C0
`define CUBE_LUT_B3E9 16'hB3C1
`define CUBE_LUT_B3EA 16'hB3C2
`define CUBE_LUT_B3EB 16'hB3C3
`define CUBE_LUT_B3EC 16'hB3C4
`define CUBE_LUT_B3ED 16'hB3C5
`define CUBE_LUT_B3EE 16'hB3C5
`define CUBE_LUT_B3EF 16'hB3C6
`define CUBE_LUT_B3F0 16'hB3C7
`define CUBE_LUT_B3F1 16'hB3C8
`define CUBE_LUT_B3F2 16'hB3C9
`define CUBE_LUT_B3F3 16'hB3CA
`define CUBE_LUT_B3F4 16'hB3CB
`define CUBE_LUT_B3F5 16'hB3CC
`define CUBE_LUT_B3F6 16'hB3CD
`define CUBE_LUT_B3F7 16'hB3CE
`define CUBE_LUT_B3F8 16'hB3CF
`define CUBE_LUT_B3F9 16'hB3D0
`define CUBE_LUT_B3FA 16'hB3D1
`define CUBE_LUT_B3FB 16'hB3D2
`define CUBE_LUT_B3FC 16'hB3D3
`define CUBE_LUT_B3FD 16'hB3D4
`define CUBE_LUT_B3FE 16'hB3D4
`define CUBE_LUT_B3FF 16'hB3D5
`define CUBE_LUT_B400 16'hB3D6
`define CUBE_LUT_B401 16'hB3D8
`define CUBE_LUT_B402 16'hB3DA
`define CUBE_LUT_B403 16'hB3DC
`define CUBE_LUT_B404 16'hB3DE
`define CUBE_LUT_B405 16'hB3E0
`define CUBE_LUT_B406 16'hB3E2
`define CUBE_LUT_B407 16'hB3E4
`define CUBE_LUT_B408 16'hB3E5
`define CUBE_LUT_B409 16'hB3E7
`define CUBE_LUT_B40A 16'hB3E9
`define CUBE_LUT_B40B 16'hB3EB
`define CUBE_LUT_B40C 16'hB3ED
`define CUBE_LUT_B40D 16'hB3EF
`define CUBE_LUT_B40E 16'hB3F1
`define CUBE_LUT_B40F 16'hB3F3
`define CUBE_LUT_B410 16'hB3F4
`define CUBE_LUT_B411 16'hB3F6
`define CUBE_LUT_B412 16'hB3F8
`define CUBE_LUT_B413 16'hB3FA
`define CUBE_LUT_B414 16'hB3FC
`define CUBE_LUT_B415 16'hB3FE
`define CUBE_LUT_B416 16'hB400
`define CUBE_LUT_B417 16'hB401
`define CUBE_LUT_B418 16'hB402
`define CUBE_LUT_B419 16'hB403
`define CUBE_LUT_B41A 16'hB404
`define CUBE_LUT_B41B 16'hB405
`define CUBE_LUT_B41C 16'hB405
`define CUBE_LUT_B41D 16'hB406
`define CUBE_LUT_B41E 16'hB407
`define CUBE_LUT_B41F 16'hB408
`define CUBE_LUT_B420 16'hB409
`define CUBE_LUT_B421 16'hB40A
`define CUBE_LUT_B422 16'hB40B
`define CUBE_LUT_B423 16'hB40C
`define CUBE_LUT_B424 16'hB40D
`define CUBE_LUT_B425 16'hB40E
`define CUBE_LUT_B426 16'hB40F
`define CUBE_LUT_B427 16'hB410
`define CUBE_LUT_B428 16'hB411
`define CUBE_LUT_B429 16'hB412
`define CUBE_LUT_B42A 16'hB413
`define CUBE_LUT_B42B 16'hB414
`define CUBE_LUT_B42C 16'hB414
`define CUBE_LUT_B42D 16'hB415
`define CUBE_LUT_B42E 16'hB416
`define CUBE_LUT_B42F 16'hB417
`define CUBE_LUT_B430 16'hB418
`define CUBE_LUT_B431 16'hB419
`define CUBE_LUT_B432 16'hB41A
`define CUBE_LUT_B433 16'hB41B
`define CUBE_LUT_B434 16'hB41C
`define CUBE_LUT_B435 16'hB41D
`define CUBE_LUT_B436 16'hB41E
`define CUBE_LUT_B437 16'hB41F
`define CUBE_LUT_B438 16'hB420
`define CUBE_LUT_B439 16'hB421
`define CUBE_LUT_B43A 16'hB422
`define CUBE_LUT_B43B 16'hB422
`define CUBE_LUT_B43C 16'hB423
`define CUBE_LUT_B43D 16'hB424
`define CUBE_LUT_B43E 16'hB425
`define CUBE_LUT_B43F 16'hB426
`define CUBE_LUT_B440 16'hB427
`define CUBE_LUT_B441 16'hB428
`define CUBE_LUT_B442 16'hB429
`define CUBE_LUT_B443 16'hB42A
`define CUBE_LUT_B444 16'hB42B
`define CUBE_LUT_B445 16'hB42C
`define CUBE_LUT_B446 16'hB42D
`define CUBE_LUT_B447 16'hB42E
`define CUBE_LUT_B448 16'hB42F
`define CUBE_LUT_B449 16'hB430
`define CUBE_LUT_B44A 16'hB430
`define CUBE_LUT_B44B 16'hB431
`define CUBE_LUT_B44C 16'hB432
`define CUBE_LUT_B44D 16'hB433
`define CUBE_LUT_B44E 16'hB434
`define CUBE_LUT_B44F 16'hB435
`define CUBE_LUT_B450 16'hB436
`define CUBE_LUT_B451 16'hB437
`define CUBE_LUT_B452 16'hB438
`define CUBE_LUT_B453 16'hB439
`define CUBE_LUT_B454 16'hB43A
`define CUBE_LUT_B455 16'hB43B
`define CUBE_LUT_B456 16'hB43C
`define CUBE_LUT_B457 16'hB43D
`define CUBE_LUT_B458 16'hB43D
`define CUBE_LUT_B459 16'hB43E
`define CUBE_LUT_B45A 16'hB43F
`define CUBE_LUT_B45B 16'hB440
`define CUBE_LUT_B45C 16'hB441
`define CUBE_LUT_B45D 16'hB442
`define CUBE_LUT_B45E 16'hB443
`define CUBE_LUT_B45F 16'hB444
`define CUBE_LUT_B460 16'hB445
`define CUBE_LUT_B461 16'hB446
`define CUBE_LUT_B462 16'hB447
`define CUBE_LUT_B463 16'hB448
`define CUBE_LUT_B464 16'hB449
`define CUBE_LUT_B465 16'hB44A
`define CUBE_LUT_B466 16'hB44A
`define CUBE_LUT_B467 16'hB44B
`define CUBE_LUT_B468 16'hB44C
`define CUBE_LUT_B469 16'hB44D
`define CUBE_LUT_B46A 16'hB44E
`define CUBE_LUT_B46B 16'hB44F
`define CUBE_LUT_B46C 16'hB450
`define CUBE_LUT_B46D 16'hB451
`define CUBE_LUT_B46E 16'hB452
`define CUBE_LUT_B46F 16'hB453
`define CUBE_LUT_B470 16'hB454
`define CUBE_LUT_B471 16'hB455
`define CUBE_LUT_B472 16'hB456
`define CUBE_LUT_B473 16'hB457
`define CUBE_LUT_B474 16'hB457
`define CUBE_LUT_B475 16'hB458
`define CUBE_LUT_B476 16'hB459
`define CUBE_LUT_B477 16'hB45A
`define CUBE_LUT_B478 16'hB45B
`define CUBE_LUT_B479 16'hB45C
`define CUBE_LUT_B47A 16'hB45D
`define CUBE_LUT_B47B 16'hB45E
`define CUBE_LUT_B47C 16'hB45F
`define CUBE_LUT_B47D 16'hB460
`define CUBE_LUT_B47E 16'hB461
`define CUBE_LUT_B47F 16'hB462
`define CUBE_LUT_B480 16'hB463
`define CUBE_LUT_B481 16'hB463
`define CUBE_LUT_B482 16'hB464
`define CUBE_LUT_B483 16'hB465
`define CUBE_LUT_B484 16'hB466
`define CUBE_LUT_B485 16'hB467
`define CUBE_LUT_B486 16'hB468
`define CUBE_LUT_B487 16'hB469
`define CUBE_LUT_B488 16'hB46A
`define CUBE_LUT_B489 16'hB46B
`define CUBE_LUT_B48A 16'hB46C
`define CUBE_LUT_B48B 16'hB46D
`define CUBE_LUT_B48C 16'hB46E
`define CUBE_LUT_B48D 16'hB46F
`define CUBE_LUT_B48E 16'hB46F
`define CUBE_LUT_B48F 16'hB470
`define CUBE_LUT_B490 16'hB471
`define CUBE_LUT_B491 16'hB472
`define CUBE_LUT_B492 16'hB473
`define CUBE_LUT_B493 16'hB474
`define CUBE_LUT_B494 16'hB475
`define CUBE_LUT_B495 16'hB476
`define CUBE_LUT_B496 16'hB477
`define CUBE_LUT_B497 16'hB478
`define CUBE_LUT_B498 16'hB479
`define CUBE_LUT_B499 16'hB47A
`define CUBE_LUT_B49A 16'hB47B
`define CUBE_LUT_B49B 16'hB47B
`define CUBE_LUT_B49C 16'hB47C
`define CUBE_LUT_B49D 16'hB47D
`define CUBE_LUT_B49E 16'hB47E
`define CUBE_LUT_B49F 16'hB47F
`define CUBE_LUT_B4A0 16'hB480
`define CUBE_LUT_B4A1 16'hB481
`define CUBE_LUT_B4A2 16'hB482
`define CUBE_LUT_B4A3 16'hB483
`define CUBE_LUT_B4A4 16'hB484
`define CUBE_LUT_B4A5 16'hB485
`define CUBE_LUT_B4A6 16'hB486
`define CUBE_LUT_B4A7 16'hB487
`define CUBE_LUT_B4A8 16'hB487
`define CUBE_LUT_B4A9 16'hB488
`define CUBE_LUT_B4AA 16'hB489
`define CUBE_LUT_B4AB 16'hB48A
`define CUBE_LUT_B4AC 16'hB48B
`define CUBE_LUT_B4AD 16'hB48C
`define CUBE_LUT_B4AE 16'hB48D
`define CUBE_LUT_B4AF 16'hB48E
`define CUBE_LUT_B4B0 16'hB48F
`define CUBE_LUT_B4B1 16'hB490
`define CUBE_LUT_B4B2 16'hB491
`define CUBE_LUT_B4B3 16'hB492
`define CUBE_LUT_B4B4 16'hB492
`define CUBE_LUT_B4B5 16'hB493
`define CUBE_LUT_B4B6 16'hB494
`define CUBE_LUT_B4B7 16'hB495
`define CUBE_LUT_B4B8 16'hB496
`define CUBE_LUT_B4B9 16'hB497
`define CUBE_LUT_B4BA 16'hB498
`define CUBE_LUT_B4BB 16'hB499
`define CUBE_LUT_B4BC 16'hB49A
`define CUBE_LUT_B4BD 16'hB49B
`define CUBE_LUT_B4BE 16'hB49C
`define CUBE_LUT_B4BF 16'hB49D
`define CUBE_LUT_B4C0 16'hB49D
`define CUBE_LUT_B4C1 16'hB49E
`define CUBE_LUT_B4C2 16'hB49F
`define CUBE_LUT_B4C3 16'hB4A0
`define CUBE_LUT_B4C4 16'hB4A1
`define CUBE_LUT_B4C5 16'hB4A2
`define CUBE_LUT_B4C6 16'hB4A3
`define CUBE_LUT_B4C7 16'hB4A4
`define CUBE_LUT_B4C8 16'hB4A5
`define CUBE_LUT_B4C9 16'hB4A6
`define CUBE_LUT_B4CA 16'hB4A7
`define CUBE_LUT_B4CB 16'hB4A8
`define CUBE_LUT_B4CC 16'hB4A8
`define CUBE_LUT_B4CD 16'hB4A9
`define CUBE_LUT_B4CE 16'hB4AA
`define CUBE_LUT_B4CF 16'hB4AB
`define CUBE_LUT_B4D0 16'hB4AC
`define CUBE_LUT_B4D1 16'hB4AD
`define CUBE_LUT_B4D2 16'hB4AE
`define CUBE_LUT_B4D3 16'hB4AF
`define CUBE_LUT_B4D4 16'hB4B0
`define CUBE_LUT_B4D5 16'hB4B1
`define CUBE_LUT_B4D6 16'hB4B2
`define CUBE_LUT_B4D7 16'hB4B3
`define CUBE_LUT_B4D8 16'hB4B3
`define CUBE_LUT_B4D9 16'hB4B4
`define CUBE_LUT_B4DA 16'hB4B5
`define CUBE_LUT_B4DB 16'hB4B6
`define CUBE_LUT_B4DC 16'hB4B7
`define CUBE_LUT_B4DD 16'hB4B8
`define CUBE_LUT_B4DE 16'hB4B9
`define CUBE_LUT_B4DF 16'hB4BA
`define CUBE_LUT_B4E0 16'hB4BB
`define CUBE_LUT_B4E1 16'hB4BC
`define CUBE_LUT_B4E2 16'hB4BD
`define CUBE_LUT_B4E3 16'hB4BE
`define CUBE_LUT_B4E4 16'hB4BE
`define CUBE_LUT_B4E5 16'hB4BF
`define CUBE_LUT_B4E6 16'hB4C0
`define CUBE_LUT_B4E7 16'hB4C1
`define CUBE_LUT_B4E8 16'hB4C2
`define CUBE_LUT_B4E9 16'hB4C3
`define CUBE_LUT_B4EA 16'hB4C4
`define CUBE_LUT_B4EB 16'hB4C5
`define CUBE_LUT_B4EC 16'hB4C6
`define CUBE_LUT_B4ED 16'hB4C7
`define CUBE_LUT_B4EE 16'hB4C8
`define CUBE_LUT_B4EF 16'hB4C8
`define CUBE_LUT_B4F0 16'hB4C9
`define CUBE_LUT_B4F1 16'hB4CA
`define CUBE_LUT_B4F2 16'hB4CB
`define CUBE_LUT_B4F3 16'hB4CC
`define CUBE_LUT_B4F4 16'hB4CD
`define CUBE_LUT_B4F5 16'hB4CE
`define CUBE_LUT_B4F6 16'hB4CF
`define CUBE_LUT_B4F7 16'hB4D0
`define CUBE_LUT_B4F8 16'hB4D1
`define CUBE_LUT_B4F9 16'hB4D2
`define CUBE_LUT_B4FA 16'hB4D2
`define CUBE_LUT_B4FB 16'hB4D3
`define CUBE_LUT_B4FC 16'hB4D4
`define CUBE_LUT_B4FD 16'hB4D5
`define CUBE_LUT_B4FE 16'hB4D6
`define CUBE_LUT_B4FF 16'hB4D7
`define CUBE_LUT_B500 16'hB4D8
`define CUBE_LUT_B501 16'hB4D9
`define CUBE_LUT_B502 16'hB4DA
`define CUBE_LUT_B503 16'hB4DB
`define CUBE_LUT_B504 16'hB4DC
`define CUBE_LUT_B505 16'hB4DC
`define CUBE_LUT_B506 16'hB4DD
`define CUBE_LUT_B507 16'hB4DE
`define CUBE_LUT_B508 16'hB4DF
`define CUBE_LUT_B509 16'hB4E0
`define CUBE_LUT_B50A 16'hB4E1
`define CUBE_LUT_B50B 16'hB4E2
`define CUBE_LUT_B50C 16'hB4E3
`define CUBE_LUT_B50D 16'hB4E4
`define CUBE_LUT_B50E 16'hB4E5
`define CUBE_LUT_B50F 16'hB4E6
`define CUBE_LUT_B510 16'hB4E6
`define CUBE_LUT_B511 16'hB4E7
`define CUBE_LUT_B512 16'hB4E8
`define CUBE_LUT_B513 16'hB4E9
`define CUBE_LUT_B514 16'hB4EA
`define CUBE_LUT_B515 16'hB4EB
`define CUBE_LUT_B516 16'hB4EC
`define CUBE_LUT_B517 16'hB4ED
`define CUBE_LUT_B518 16'hB4EE
`define CUBE_LUT_B519 16'hB4EF
`define CUBE_LUT_B51A 16'hB4EF
`define CUBE_LUT_B51B 16'hB4F0
`define CUBE_LUT_B51C 16'hB4F1
`define CUBE_LUT_B51D 16'hB4F2
`define CUBE_LUT_B51E 16'hB4F3
`define CUBE_LUT_B51F 16'hB4F4
`define CUBE_LUT_B520 16'hB4F5
`define CUBE_LUT_B521 16'hB4F6
`define CUBE_LUT_B522 16'hB4F7
`define CUBE_LUT_B523 16'hB4F8
`define CUBE_LUT_B524 16'hB4F9
`define CUBE_LUT_B525 16'hB4F9
`define CUBE_LUT_B526 16'hB4FA
`define CUBE_LUT_B527 16'hB4FB
`define CUBE_LUT_B528 16'hB4FC
`define CUBE_LUT_B529 16'hB4FD
`define CUBE_LUT_B52A 16'hB4FE
`define CUBE_LUT_B52B 16'hB4FF
`define CUBE_LUT_B52C 16'hB500
`define CUBE_LUT_B52D 16'hB501
`define CUBE_LUT_B52E 16'hB502
`define CUBE_LUT_B52F 16'hB502
`define CUBE_LUT_B530 16'hB503
`define CUBE_LUT_B531 16'hB504
`define CUBE_LUT_B532 16'hB505
`define CUBE_LUT_B533 16'hB506
`define CUBE_LUT_B534 16'hB507
`define CUBE_LUT_B535 16'hB508
`define CUBE_LUT_B536 16'hB509
`define CUBE_LUT_B537 16'hB50A
`define CUBE_LUT_B538 16'hB50B
`define CUBE_LUT_B539 16'hB50B
`define CUBE_LUT_B53A 16'hB50C
`define CUBE_LUT_B53B 16'hB50D
`define CUBE_LUT_B53C 16'hB50E
`define CUBE_LUT_B53D 16'hB50F
`define CUBE_LUT_B53E 16'hB510
`define CUBE_LUT_B53F 16'hB511
`define CUBE_LUT_B540 16'hB512
`define CUBE_LUT_B541 16'hB513
`define CUBE_LUT_B542 16'hB514
`define CUBE_LUT_B543 16'hB514
`define CUBE_LUT_B544 16'hB515
`define CUBE_LUT_B545 16'hB516
`define CUBE_LUT_B546 16'hB517
`define CUBE_LUT_B547 16'hB518
`define CUBE_LUT_B548 16'hB519
`define CUBE_LUT_B549 16'hB51A
`define CUBE_LUT_B54A 16'hB51B
`define CUBE_LUT_B54B 16'hB51C
`define CUBE_LUT_B54C 16'hB51D
`define CUBE_LUT_B54D 16'hB51D
`define CUBE_LUT_B54E 16'hB51E
`define CUBE_LUT_B54F 16'hB51F
`define CUBE_LUT_B550 16'hB520
`define CUBE_LUT_B551 16'hB521
`define CUBE_LUT_B552 16'hB522
`define CUBE_LUT_B553 16'hB523
`define CUBE_LUT_B554 16'hB524
`define CUBE_LUT_B555 16'hB525
`define CUBE_LUT_B556 16'hB526
`define CUBE_LUT_B557 16'hB526
`define CUBE_LUT_B558 16'hB527
`define CUBE_LUT_B559 16'hB528
`define CUBE_LUT_B55A 16'hB529
`define CUBE_LUT_B55B 16'hB52A
`define CUBE_LUT_B55C 16'hB52B
`define CUBE_LUT_B55D 16'hB52C
`define CUBE_LUT_B55E 16'hB52D
`define CUBE_LUT_B55F 16'hB52E
`define CUBE_LUT_B560 16'hB52E
`define CUBE_LUT_B561 16'hB52F
`define CUBE_LUT_B562 16'hB530
`define CUBE_LUT_B563 16'hB531
`define CUBE_LUT_B564 16'hB532
`define CUBE_LUT_B565 16'hB533
`define CUBE_LUT_B566 16'hB534
`define CUBE_LUT_B567 16'hB535
`define CUBE_LUT_B568 16'hB536
`define CUBE_LUT_B569 16'hB537
`define CUBE_LUT_B56A 16'hB537
`define CUBE_LUT_B56B 16'hB538
`define CUBE_LUT_B56C 16'hB539
`define CUBE_LUT_B56D 16'hB53A
`define CUBE_LUT_B56E 16'hB53B
`define CUBE_LUT_B56F 16'hB53C
`define CUBE_LUT_B570 16'hB53D
`define CUBE_LUT_B571 16'hB53E
`define CUBE_LUT_B572 16'hB53F
`define CUBE_LUT_B573 16'hB53F
`define CUBE_LUT_B574 16'hB540
`define CUBE_LUT_B575 16'hB541
`define CUBE_LUT_B576 16'hB542
`define CUBE_LUT_B577 16'hB543
`define CUBE_LUT_B578 16'hB544
`define CUBE_LUT_B579 16'hB545
`define CUBE_LUT_B57A 16'hB546
`define CUBE_LUT_B57B 16'hB547
`define CUBE_LUT_B57C 16'hB547
`define CUBE_LUT_B57D 16'hB548
`define CUBE_LUT_B57E 16'hB549
`define CUBE_LUT_B57F 16'hB54A
`define CUBE_LUT_B580 16'hB54B
`define CUBE_LUT_B581 16'hB54C
`define CUBE_LUT_B582 16'hB54D
`define CUBE_LUT_B583 16'hB54E
`define CUBE_LUT_B584 16'hB54F
`define CUBE_LUT_B585 16'hB54F
`define CUBE_LUT_B586 16'hB550
`define CUBE_LUT_B587 16'hB551
`define CUBE_LUT_B588 16'hB552
`define CUBE_LUT_B589 16'hB553
`define CUBE_LUT_B58A 16'hB554
`define CUBE_LUT_B58B 16'hB555
`define CUBE_LUT_B58C 16'hB556
`define CUBE_LUT_B58D 16'hB557
`define CUBE_LUT_B58E 16'hB557
`define CUBE_LUT_B58F 16'hB558
`define CUBE_LUT_B590 16'hB559
`define CUBE_LUT_B591 16'hB55A
`define CUBE_LUT_B592 16'hB55B
`define CUBE_LUT_B593 16'hB55C
`define CUBE_LUT_B594 16'hB55D
`define CUBE_LUT_B595 16'hB55E
`define CUBE_LUT_B596 16'hB55F
`define CUBE_LUT_B597 16'hB55F
`define CUBE_LUT_B598 16'hB560
`define CUBE_LUT_B599 16'hB561
`define CUBE_LUT_B59A 16'hB562
`define CUBE_LUT_B59B 16'hB563
`define CUBE_LUT_B59C 16'hB564
`define CUBE_LUT_B59D 16'hB565
`define CUBE_LUT_B59E 16'hB566
`define CUBE_LUT_B59F 16'hB567
`define CUBE_LUT_B5A0 16'hB567
`define CUBE_LUT_B5A1 16'hB568
`define CUBE_LUT_B5A2 16'hB569
`define CUBE_LUT_B5A3 16'hB56A
`define CUBE_LUT_B5A4 16'hB56B
`define CUBE_LUT_B5A5 16'hB56C
`define CUBE_LUT_B5A6 16'hB56D
`define CUBE_LUT_B5A7 16'hB56E
`define CUBE_LUT_B5A8 16'hB56F
`define CUBE_LUT_B5A9 16'hB56F
`define CUBE_LUT_B5AA 16'hB570
`define CUBE_LUT_B5AB 16'hB571
`define CUBE_LUT_B5AC 16'hB572
`define CUBE_LUT_B5AD 16'hB573
`define CUBE_LUT_B5AE 16'hB574
`define CUBE_LUT_B5AF 16'hB575
`define CUBE_LUT_B5B0 16'hB576
`define CUBE_LUT_B5B1 16'hB577
`define CUBE_LUT_B5B2 16'hB577
`define CUBE_LUT_B5B3 16'hB578
`define CUBE_LUT_B5B4 16'hB579
`define CUBE_LUT_B5B5 16'hB57A
`define CUBE_LUT_B5B6 16'hB57B
`define CUBE_LUT_B5B7 16'hB57C
`define CUBE_LUT_B5B8 16'hB57D
`define CUBE_LUT_B5B9 16'hB57E
`define CUBE_LUT_B5BA 16'hB57E
`define CUBE_LUT_B5BB 16'hB57F
`define CUBE_LUT_B5BC 16'hB580
`define CUBE_LUT_B5BD 16'hB581
`define CUBE_LUT_B5BE 16'hB582
`define CUBE_LUT_B5BF 16'hB583
`define CUBE_LUT_B5C0 16'hB584
`define CUBE_LUT_B5C1 16'hB585
`define CUBE_LUT_B5C2 16'hB586
`define CUBE_LUT_B5C3 16'hB586
`define CUBE_LUT_B5C4 16'hB587
`define CUBE_LUT_B5C5 16'hB588
`define CUBE_LUT_B5C6 16'hB589
`define CUBE_LUT_B5C7 16'hB58A
`define CUBE_LUT_B5C8 16'hB58B
`define CUBE_LUT_B5C9 16'hB58C
`define CUBE_LUT_B5CA 16'hB58D
`define CUBE_LUT_B5CB 16'hB58D
`define CUBE_LUT_B5CC 16'hB58E
`define CUBE_LUT_B5CD 16'hB58F
`define CUBE_LUT_B5CE 16'hB590
`define CUBE_LUT_B5CF 16'hB591
`define CUBE_LUT_B5D0 16'hB592
`define CUBE_LUT_B5D1 16'hB593
`define CUBE_LUT_B5D2 16'hB594
`define CUBE_LUT_B5D3 16'hB594
`define CUBE_LUT_B5D4 16'hB595
`define CUBE_LUT_B5D5 16'hB596
`define CUBE_LUT_B5D6 16'hB597
`define CUBE_LUT_B5D7 16'hB598
`define CUBE_LUT_B5D8 16'hB599
`define CUBE_LUT_B5D9 16'hB59A
`define CUBE_LUT_B5DA 16'hB59B
`define CUBE_LUT_B5DB 16'hB59B
`define CUBE_LUT_B5DC 16'hB59C
`define CUBE_LUT_B5DD 16'hB59D
`define CUBE_LUT_B5DE 16'hB59E
`define CUBE_LUT_B5DF 16'hB59F
`define CUBE_LUT_B5E0 16'hB5A0
`define CUBE_LUT_B5E1 16'hB5A1
`define CUBE_LUT_B5E2 16'hB5A2
`define CUBE_LUT_B5E3 16'hB5A2
`define CUBE_LUT_B5E4 16'hB5A3
`define CUBE_LUT_B5E5 16'hB5A4
`define CUBE_LUT_B5E6 16'hB5A5
`define CUBE_LUT_B5E7 16'hB5A6
`define CUBE_LUT_B5E8 16'hB5A7
`define CUBE_LUT_B5E9 16'hB5A8
`define CUBE_LUT_B5EA 16'hB5A9
`define CUBE_LUT_B5EB 16'hB5A9
`define CUBE_LUT_B5EC 16'hB5AA
`define CUBE_LUT_B5ED 16'hB5AB
`define CUBE_LUT_B5EE 16'hB5AC
`define CUBE_LUT_B5EF 16'hB5AD
`define CUBE_LUT_B5F0 16'hB5AE
`define CUBE_LUT_B5F1 16'hB5AF
`define CUBE_LUT_B5F2 16'hB5B0
`define CUBE_LUT_B5F3 16'hB5B0
`define CUBE_LUT_B5F4 16'hB5B1
`define CUBE_LUT_B5F5 16'hB5B2
`define CUBE_LUT_B5F6 16'hB5B3
`define CUBE_LUT_B5F7 16'hB5B4
`define CUBE_LUT_B5F8 16'hB5B5
`define CUBE_LUT_B5F9 16'hB5B6
`define CUBE_LUT_B5FA 16'hB5B7
`define CUBE_LUT_B5FB 16'hB5B7
`define CUBE_LUT_B5FC 16'hB5B8
`define CUBE_LUT_B5FD 16'hB5B9
`define CUBE_LUT_B5FE 16'hB5BA
`define CUBE_LUT_B5FF 16'hB5BB
`define CUBE_LUT_B600 16'hB5BC
`define CUBE_LUT_B601 16'hB5BD
`define CUBE_LUT_B602 16'hB5BE
`define CUBE_LUT_B603 16'hB5BE
`define CUBE_LUT_B604 16'hB5BF
`define CUBE_LUT_B605 16'hB5C0
`define CUBE_LUT_B606 16'hB5C1
`define CUBE_LUT_B607 16'hB5C2
`define CUBE_LUT_B608 16'hB5C3
`define CUBE_LUT_B609 16'hB5C4
`define CUBE_LUT_B60A 16'hB5C5
`define CUBE_LUT_B60B 16'hB5C5
`define CUBE_LUT_B60C 16'hB5C6
`define CUBE_LUT_B60D 16'hB5C7
`define CUBE_LUT_B60E 16'hB5C8
`define CUBE_LUT_B60F 16'hB5C9
`define CUBE_LUT_B610 16'hB5CA
`define CUBE_LUT_B611 16'hB5CB
`define CUBE_LUT_B612 16'hB5CB
`define CUBE_LUT_B613 16'hB5CC
`define CUBE_LUT_B614 16'hB5CD
`define CUBE_LUT_B615 16'hB5CE
`define CUBE_LUT_B616 16'hB5CF
`define CUBE_LUT_B617 16'hB5D0
`define CUBE_LUT_B618 16'hB5D1
`define CUBE_LUT_B619 16'hB5D2
`define CUBE_LUT_B61A 16'hB5D2
`define CUBE_LUT_B61B 16'hB5D3
`define CUBE_LUT_B61C 16'hB5D4
`define CUBE_LUT_B61D 16'hB5D5
`define CUBE_LUT_B61E 16'hB5D6
`define CUBE_LUT_B61F 16'hB5D7
`define CUBE_LUT_B620 16'hB5D8
`define CUBE_LUT_B621 16'hB5D9
`define CUBE_LUT_B622 16'hB5D9
`define CUBE_LUT_B623 16'hB5DA
`define CUBE_LUT_B624 16'hB5DB
`define CUBE_LUT_B625 16'hB5DC
`define CUBE_LUT_B626 16'hB5DD
`define CUBE_LUT_B627 16'hB5DE
`define CUBE_LUT_B628 16'hB5DF
`define CUBE_LUT_B629 16'hB5DF
`define CUBE_LUT_B62A 16'hB5E0
`define CUBE_LUT_B62B 16'hB5E1
`define CUBE_LUT_B62C 16'hB5E2
`define CUBE_LUT_B62D 16'hB5E3
`define CUBE_LUT_B62E 16'hB5E4
`define CUBE_LUT_B62F 16'hB5E5
`define CUBE_LUT_B630 16'hB5E5
`define CUBE_LUT_B631 16'hB5E6
`define CUBE_LUT_B632 16'hB5E7
`define CUBE_LUT_B633 16'hB5E8
`define CUBE_LUT_B634 16'hB5E9
`define CUBE_LUT_B635 16'hB5EA
`define CUBE_LUT_B636 16'hB5EB
`define CUBE_LUT_B637 16'hB5EC
`define CUBE_LUT_B638 16'hB5EC
`define CUBE_LUT_B639 16'hB5ED
`define CUBE_LUT_B63A 16'hB5EE
`define CUBE_LUT_B63B 16'hB5EF
`define CUBE_LUT_B63C 16'hB5F0
`define CUBE_LUT_B63D 16'hB5F1
`define CUBE_LUT_B63E 16'hB5F2
`define CUBE_LUT_B63F 16'hB5F2
`define CUBE_LUT_B640 16'hB5F3
`define CUBE_LUT_B641 16'hB5F4
`define CUBE_LUT_B642 16'hB5F5
`define CUBE_LUT_B643 16'hB5F6
`define CUBE_LUT_B644 16'hB5F7
`define CUBE_LUT_B645 16'hB5F8
`define CUBE_LUT_B646 16'hB5F8
`define CUBE_LUT_B647 16'hB5F9
`define CUBE_LUT_B648 16'hB5FA
`define CUBE_LUT_B649 16'hB5FB
`define CUBE_LUT_B64A 16'hB5FC
`define CUBE_LUT_B64B 16'hB5FD
`define CUBE_LUT_B64C 16'hB5FE
`define CUBE_LUT_B64D 16'hB5FE
`define CUBE_LUT_B64E 16'hB5FF
`define CUBE_LUT_B64F 16'hB600
`define CUBE_LUT_B650 16'hB601
`define CUBE_LUT_B651 16'hB602
`define CUBE_LUT_B652 16'hB603
`define CUBE_LUT_B653 16'hB604
`define CUBE_LUT_B654 16'hB605
`define CUBE_LUT_B655 16'hB605
`define CUBE_LUT_B656 16'hB606
`define CUBE_LUT_B657 16'hB607
`define CUBE_LUT_B658 16'hB608
`define CUBE_LUT_B659 16'hB609
`define CUBE_LUT_B65A 16'hB60A
`define CUBE_LUT_B65B 16'hB60B
`define CUBE_LUT_B65C 16'hB60B
`define CUBE_LUT_B65D 16'hB60C
`define CUBE_LUT_B65E 16'hB60D
`define CUBE_LUT_B65F 16'hB60E
`define CUBE_LUT_B660 16'hB60F
`define CUBE_LUT_B661 16'hB610
`define CUBE_LUT_B662 16'hB611
`define CUBE_LUT_B663 16'hB611
`define CUBE_LUT_B664 16'hB612
`define CUBE_LUT_B665 16'hB613
`define CUBE_LUT_B666 16'hB614
`define CUBE_LUT_B667 16'hB615
`define CUBE_LUT_B668 16'hB616
`define CUBE_LUT_B669 16'hB616
`define CUBE_LUT_B66A 16'hB617
`define CUBE_LUT_B66B 16'hB618
`define CUBE_LUT_B66C 16'hB619
`define CUBE_LUT_B66D 16'hB61A
`define CUBE_LUT_B66E 16'hB61B
`define CUBE_LUT_B66F 16'hB61C
`define CUBE_LUT_B670 16'hB61C
`define CUBE_LUT_B671 16'hB61D
`define CUBE_LUT_B672 16'hB61E
`define CUBE_LUT_B673 16'hB61F
`define CUBE_LUT_B674 16'hB620
`define CUBE_LUT_B675 16'hB621
`define CUBE_LUT_B676 16'hB622
`define CUBE_LUT_B677 16'hB622
`define CUBE_LUT_B678 16'hB623
`define CUBE_LUT_B679 16'hB624
`define CUBE_LUT_B67A 16'hB625
`define CUBE_LUT_B67B 16'hB626
`define CUBE_LUT_B67C 16'hB627
`define CUBE_LUT_B67D 16'hB628
`define CUBE_LUT_B67E 16'hB628
`define CUBE_LUT_B67F 16'hB629
`define CUBE_LUT_B680 16'hB62A
`define CUBE_LUT_B681 16'hB62B
`define CUBE_LUT_B682 16'hB62C
`define CUBE_LUT_B683 16'hB62D
`define CUBE_LUT_B684 16'hB62E
`define CUBE_LUT_B685 16'hB62E
`define CUBE_LUT_B686 16'hB62F
`define CUBE_LUT_B687 16'hB630
`define CUBE_LUT_B688 16'hB631
`define CUBE_LUT_B689 16'hB632
`define CUBE_LUT_B68A 16'hB633
`define CUBE_LUT_B68B 16'hB633
`define CUBE_LUT_B68C 16'hB634
`define CUBE_LUT_B68D 16'hB635
`define CUBE_LUT_B68E 16'hB636
`define CUBE_LUT_B68F 16'hB637
`define CUBE_LUT_B690 16'hB638
`define CUBE_LUT_B691 16'hB639
`define CUBE_LUT_B692 16'hB639
`define CUBE_LUT_B693 16'hB63A
`define CUBE_LUT_B694 16'hB63B
`define CUBE_LUT_B695 16'hB63C
`define CUBE_LUT_B696 16'hB63D
`define CUBE_LUT_B697 16'hB63E
`define CUBE_LUT_B698 16'hB63F
`define CUBE_LUT_B699 16'hB63F
`define CUBE_LUT_B69A 16'hB640
`define CUBE_LUT_B69B 16'hB641
`define CUBE_LUT_B69C 16'hB642
`define CUBE_LUT_B69D 16'hB643
`define CUBE_LUT_B69E 16'hB644
`define CUBE_LUT_B69F 16'hB644
`define CUBE_LUT_B6A0 16'hB645
`define CUBE_LUT_B6A1 16'hB646
`define CUBE_LUT_B6A2 16'hB647
`define CUBE_LUT_B6A3 16'hB648
`define CUBE_LUT_B6A4 16'hB649
`define CUBE_LUT_B6A5 16'hB64A
`define CUBE_LUT_B6A6 16'hB64A
`define CUBE_LUT_B6A7 16'hB64B
`define CUBE_LUT_B6A8 16'hB64C
`define CUBE_LUT_B6A9 16'hB64D
`define CUBE_LUT_B6AA 16'hB64E
`define CUBE_LUT_B6AB 16'hB64F
`define CUBE_LUT_B6AC 16'hB64F
`define CUBE_LUT_B6AD 16'hB650
`define CUBE_LUT_B6AE 16'hB651
`define CUBE_LUT_B6AF 16'hB652
`define CUBE_LUT_B6B0 16'hB653
`define CUBE_LUT_B6B1 16'hB654
`define CUBE_LUT_B6B2 16'hB654
`define CUBE_LUT_B6B3 16'hB655
`define CUBE_LUT_B6B4 16'hB656
`define CUBE_LUT_B6B5 16'hB657
`define CUBE_LUT_B6B6 16'hB658
`define CUBE_LUT_B6B7 16'hB659
`define CUBE_LUT_B6B8 16'hB65A
`define CUBE_LUT_B6B9 16'hB65A
`define CUBE_LUT_B6BA 16'hB65B
`define CUBE_LUT_B6BB 16'hB65C
`define CUBE_LUT_B6BC 16'hB65D
`define CUBE_LUT_B6BD 16'hB65E
`define CUBE_LUT_B6BE 16'hB65F
`define CUBE_LUT_B6BF 16'hB65F
`define CUBE_LUT_B6C0 16'hB660
`define CUBE_LUT_B6C1 16'hB661
`define CUBE_LUT_B6C2 16'hB662
`define CUBE_LUT_B6C3 16'hB663
`define CUBE_LUT_B6C4 16'hB664
`define CUBE_LUT_B6C5 16'hB664
`define CUBE_LUT_B6C6 16'hB665
`define CUBE_LUT_B6C7 16'hB666
`define CUBE_LUT_B6C8 16'hB667
`define CUBE_LUT_B6C9 16'hB668
`define CUBE_LUT_B6CA 16'hB669
`define CUBE_LUT_B6CB 16'hB66A
`define CUBE_LUT_B6CC 16'hB66A
`define CUBE_LUT_B6CD 16'hB66B
`define CUBE_LUT_B6CE 16'hB66C
`define CUBE_LUT_B6CF 16'hB66D
`define CUBE_LUT_B6D0 16'hB66E
`define CUBE_LUT_B6D1 16'hB66F
`define CUBE_LUT_B6D2 16'hB66F
`define CUBE_LUT_B6D3 16'hB670
`define CUBE_LUT_B6D4 16'hB671
`define CUBE_LUT_B6D5 16'hB672
`define CUBE_LUT_B6D6 16'hB673
`define CUBE_LUT_B6D7 16'hB674
`define CUBE_LUT_B6D8 16'hB674
`define CUBE_LUT_B6D9 16'hB675
`define CUBE_LUT_B6DA 16'hB676
`define CUBE_LUT_B6DB 16'hB677
`define CUBE_LUT_B6DC 16'hB678
`define CUBE_LUT_B6DD 16'hB679
`define CUBE_LUT_B6DE 16'hB679
`define CUBE_LUT_B6DF 16'hB67A
`define CUBE_LUT_B6E0 16'hB67B
`define CUBE_LUT_B6E1 16'hB67C
`define CUBE_LUT_B6E2 16'hB67D
`define CUBE_LUT_B6E3 16'hB67E
`define CUBE_LUT_B6E4 16'hB67E
`define CUBE_LUT_B6E5 16'hB67F
`define CUBE_LUT_B6E6 16'hB680
`define CUBE_LUT_B6E7 16'hB681
`define CUBE_LUT_B6E8 16'hB682
`define CUBE_LUT_B6E9 16'hB683
`define CUBE_LUT_B6EA 16'hB683
`define CUBE_LUT_B6EB 16'hB684
`define CUBE_LUT_B6EC 16'hB685
`define CUBE_LUT_B6ED 16'hB686
`define CUBE_LUT_B6EE 16'hB687
`define CUBE_LUT_B6EF 16'hB688
`define CUBE_LUT_B6F0 16'hB688
`define CUBE_LUT_B6F1 16'hB689
`define CUBE_LUT_B6F2 16'hB68A
`define CUBE_LUT_B6F3 16'hB68B
`define CUBE_LUT_B6F4 16'hB68C
`define CUBE_LUT_B6F5 16'hB68D
`define CUBE_LUT_B6F6 16'hB68D
`define CUBE_LUT_B6F7 16'hB68E
`define CUBE_LUT_B6F8 16'hB68F
`define CUBE_LUT_B6F9 16'hB690
`define CUBE_LUT_B6FA 16'hB691
`define CUBE_LUT_B6FB 16'hB692
`define CUBE_LUT_B6FC 16'hB692
`define CUBE_LUT_B6FD 16'hB693
`define CUBE_LUT_B6FE 16'hB694
`define CUBE_LUT_B6FF 16'hB695
`define CUBE_LUT_B700 16'hB696
`define CUBE_LUT_B701 16'hB697
`define CUBE_LUT_B702 16'hB697
`define CUBE_LUT_B703 16'hB698
`define CUBE_LUT_B704 16'hB699
`define CUBE_LUT_B705 16'hB69A
`define CUBE_LUT_B706 16'hB69B
`define CUBE_LUT_B707 16'hB69C
`define CUBE_LUT_B708 16'hB69C
`define CUBE_LUT_B709 16'hB69D
`define CUBE_LUT_B70A 16'hB69E
`define CUBE_LUT_B70B 16'hB69F
`define CUBE_LUT_B70C 16'hB6A0
`define CUBE_LUT_B70D 16'hB6A1
`define CUBE_LUT_B70E 16'hB6A1
`define CUBE_LUT_B70F 16'hB6A2
`define CUBE_LUT_B710 16'hB6A3
`define CUBE_LUT_B711 16'hB6A4
`define CUBE_LUT_B712 16'hB6A5
`define CUBE_LUT_B713 16'hB6A6
`define CUBE_LUT_B714 16'hB6A6
`define CUBE_LUT_B715 16'hB6A7
`define CUBE_LUT_B716 16'hB6A8
`define CUBE_LUT_B717 16'hB6A9
`define CUBE_LUT_B718 16'hB6AA
`define CUBE_LUT_B719 16'hB6AB
`define CUBE_LUT_B71A 16'hB6AB
`define CUBE_LUT_B71B 16'hB6AC
`define CUBE_LUT_B71C 16'hB6AD
`define CUBE_LUT_B71D 16'hB6AE
`define CUBE_LUT_B71E 16'hB6AF
`define CUBE_LUT_B71F 16'hB6AF
`define CUBE_LUT_B720 16'hB6B0
`define CUBE_LUT_B721 16'hB6B1
`define CUBE_LUT_B722 16'hB6B2
`define CUBE_LUT_B723 16'hB6B3
`define CUBE_LUT_B724 16'hB6B4
`define CUBE_LUT_B725 16'hB6B4
`define CUBE_LUT_B726 16'hB6B5
`define CUBE_LUT_B727 16'hB6B6
`define CUBE_LUT_B728 16'hB6B7
`define CUBE_LUT_B729 16'hB6B8
`define CUBE_LUT_B72A 16'hB6B9
`define CUBE_LUT_B72B 16'hB6B9
`define CUBE_LUT_B72C 16'hB6BA
`define CUBE_LUT_B72D 16'hB6BB
`define CUBE_LUT_B72E 16'hB6BC
`define CUBE_LUT_B72F 16'hB6BD
`define CUBE_LUT_B730 16'hB6BD
`define CUBE_LUT_B731 16'hB6BE
`define CUBE_LUT_B732 16'hB6BF
`define CUBE_LUT_B733 16'hB6C0
`define CUBE_LUT_B734 16'hB6C1
`define CUBE_LUT_B735 16'hB6C2
`define CUBE_LUT_B736 16'hB6C2
`define CUBE_LUT_B737 16'hB6C3
`define CUBE_LUT_B738 16'hB6C4
`define CUBE_LUT_B739 16'hB6C5
`define CUBE_LUT_B73A 16'hB6C6
`define CUBE_LUT_B73B 16'hB6C7
`define CUBE_LUT_B73C 16'hB6C7
`define CUBE_LUT_B73D 16'hB6C8
`define CUBE_LUT_B73E 16'hB6C9
`define CUBE_LUT_B73F 16'hB6CA
`define CUBE_LUT_B740 16'hB6CB
`define CUBE_LUT_B741 16'hB6CB
`define CUBE_LUT_B742 16'hB6CC
`define CUBE_LUT_B743 16'hB6CD
`define CUBE_LUT_B744 16'hB6CE
`define CUBE_LUT_B745 16'hB6CF
`define CUBE_LUT_B746 16'hB6D0
`define CUBE_LUT_B747 16'hB6D0
`define CUBE_LUT_B748 16'hB6D1
`define CUBE_LUT_B749 16'hB6D2
`define CUBE_LUT_B74A 16'hB6D3
`define CUBE_LUT_B74B 16'hB6D4
`define CUBE_LUT_B74C 16'hB6D4
`define CUBE_LUT_B74D 16'hB6D5
`define CUBE_LUT_B74E 16'hB6D6
`define CUBE_LUT_B74F 16'hB6D7
`define CUBE_LUT_B750 16'hB6D8
`define CUBE_LUT_B751 16'hB6D9
`define CUBE_LUT_B752 16'hB6D9
`define CUBE_LUT_B753 16'hB6DA
`define CUBE_LUT_B754 16'hB6DB
`define CUBE_LUT_B755 16'hB6DC
`define CUBE_LUT_B756 16'hB6DD
`define CUBE_LUT_B757 16'hB6DD
`define CUBE_LUT_B758 16'hB6DE
`define CUBE_LUT_B759 16'hB6DF
`define CUBE_LUT_B75A 16'hB6E0
`define CUBE_LUT_B75B 16'hB6E1
`define CUBE_LUT_B75C 16'hB6E1
`define CUBE_LUT_B75D 16'hB6E2
`define CUBE_LUT_B75E 16'hB6E3
`define CUBE_LUT_B75F 16'hB6E4
`define CUBE_LUT_B760 16'hB6E5
`define CUBE_LUT_B761 16'hB6E6
`define CUBE_LUT_B762 16'hB6E6
`define CUBE_LUT_B763 16'hB6E7
`define CUBE_LUT_B764 16'hB6E8
`define CUBE_LUT_B765 16'hB6E9
`define CUBE_LUT_B766 16'hB6EA
`define CUBE_LUT_B767 16'hB6EA
`define CUBE_LUT_B768 16'hB6EB
`define CUBE_LUT_B769 16'hB6EC
`define CUBE_LUT_B76A 16'hB6ED
`define CUBE_LUT_B76B 16'hB6EE
`define CUBE_LUT_B76C 16'hB6EF
`define CUBE_LUT_B76D 16'hB6EF
`define CUBE_LUT_B76E 16'hB6F0
`define CUBE_LUT_B76F 16'hB6F1
`define CUBE_LUT_B770 16'hB6F2
`define CUBE_LUT_B771 16'hB6F3
`define CUBE_LUT_B772 16'hB6F3
`define CUBE_LUT_B773 16'hB6F4
`define CUBE_LUT_B774 16'hB6F5
`define CUBE_LUT_B775 16'hB6F6
`define CUBE_LUT_B776 16'hB6F7
`define CUBE_LUT_B777 16'hB6F7
`define CUBE_LUT_B778 16'hB6F8
`define CUBE_LUT_B779 16'hB6F9
`define CUBE_LUT_B77A 16'hB6FA
`define CUBE_LUT_B77B 16'hB6FB
`define CUBE_LUT_B77C 16'hB6FB
`define CUBE_LUT_B77D 16'hB6FC
`define CUBE_LUT_B77E 16'hB6FD
`define CUBE_LUT_B77F 16'hB6FE
`define CUBE_LUT_B780 16'hB6FF
`define CUBE_LUT_B781 16'hB700
`define CUBE_LUT_B782 16'hB700
`define CUBE_LUT_B783 16'hB701
`define CUBE_LUT_B784 16'hB702
`define CUBE_LUT_B785 16'hB703
`define CUBE_LUT_B786 16'hB704
`define CUBE_LUT_B787 16'hB704
`define CUBE_LUT_B788 16'hB705
`define CUBE_LUT_B789 16'hB706
`define CUBE_LUT_B78A 16'hB707
`define CUBE_LUT_B78B 16'hB708
`define CUBE_LUT_B78C 16'hB708
`define CUBE_LUT_B78D 16'hB709
`define CUBE_LUT_B78E 16'hB70A
`define CUBE_LUT_B78F 16'hB70B
`define CUBE_LUT_B790 16'hB70C
`define CUBE_LUT_B791 16'hB70C
`define CUBE_LUT_B792 16'hB70D
`define CUBE_LUT_B793 16'hB70E
`define CUBE_LUT_B794 16'hB70F
`define CUBE_LUT_B795 16'hB710
`define CUBE_LUT_B796 16'hB710
`define CUBE_LUT_B797 16'hB711
`define CUBE_LUT_B798 16'hB712
`define CUBE_LUT_B799 16'hB713
`define CUBE_LUT_B79A 16'hB714
`define CUBE_LUT_B79B 16'hB715
`define CUBE_LUT_B79C 16'hB715
`define CUBE_LUT_B79D 16'hB716
`define CUBE_LUT_B79E 16'hB717
`define CUBE_LUT_B79F 16'hB718
`define CUBE_LUT_B7A0 16'hB719
`define CUBE_LUT_B7A1 16'hB719
`define CUBE_LUT_B7A2 16'hB71A
`define CUBE_LUT_B7A3 16'hB71B
`define CUBE_LUT_B7A4 16'hB71C
`define CUBE_LUT_B7A5 16'hB71D
`define CUBE_LUT_B7A6 16'hB71D
`define CUBE_LUT_B7A7 16'hB71E
`define CUBE_LUT_B7A8 16'hB71F
`define CUBE_LUT_B7A9 16'hB720
`define CUBE_LUT_B7AA 16'hB721
`define CUBE_LUT_B7AB 16'hB721
`define CUBE_LUT_B7AC 16'hB722
`define CUBE_LUT_B7AD 16'hB723
`define CUBE_LUT_B7AE 16'hB724
`define CUBE_LUT_B7AF 16'hB725
`define CUBE_LUT_B7B0 16'hB725
`define CUBE_LUT_B7B1 16'hB726
`define CUBE_LUT_B7B2 16'hB727
`define CUBE_LUT_B7B3 16'hB728
`define CUBE_LUT_B7B4 16'hB729
`define CUBE_LUT_B7B5 16'hB729
`define CUBE_LUT_B7B6 16'hB72A
`define CUBE_LUT_B7B7 16'hB72B
`define CUBE_LUT_B7B8 16'hB72C
`define CUBE_LUT_B7B9 16'hB72D
`define CUBE_LUT_B7BA 16'hB72D
`define CUBE_LUT_B7BB 16'hB72E
`define CUBE_LUT_B7BC 16'hB72F
`define CUBE_LUT_B7BD 16'hB730
`define CUBE_LUT_B7BE 16'hB731
`define CUBE_LUT_B7BF 16'hB731
`define CUBE_LUT_B7C0 16'hB732
`define CUBE_LUT_B7C1 16'hB733
`define CUBE_LUT_B7C2 16'hB734
`define CUBE_LUT_B7C3 16'hB735
`define CUBE_LUT_B7C4 16'hB735
`define CUBE_LUT_B7C5 16'hB736
`define CUBE_LUT_B7C6 16'hB737
`define CUBE_LUT_B7C7 16'hB738
`define CUBE_LUT_B7C8 16'hB739
`define CUBE_LUT_B7C9 16'hB739
`define CUBE_LUT_B7CA 16'hB73A
`define CUBE_LUT_B7CB 16'hB73B
`define CUBE_LUT_B7CC 16'hB73C
`define CUBE_LUT_B7CD 16'hB73C
`define CUBE_LUT_B7CE 16'hB73D
`define CUBE_LUT_B7CF 16'hB73E
`define CUBE_LUT_B7D0 16'hB73F
`define CUBE_LUT_B7D1 16'hB740
`define CUBE_LUT_B7D2 16'hB740
`define CUBE_LUT_B7D3 16'hB741
`define CUBE_LUT_B7D4 16'hB742
`define CUBE_LUT_B7D5 16'hB743
`define CUBE_LUT_B7D6 16'hB744
`define CUBE_LUT_B7D7 16'hB744
`define CUBE_LUT_B7D8 16'hB745
`define CUBE_LUT_B7D9 16'hB746
`define CUBE_LUT_B7DA 16'hB747
`define CUBE_LUT_B7DB 16'hB748
`define CUBE_LUT_B7DC 16'hB748
`define CUBE_LUT_B7DD 16'hB749
`define CUBE_LUT_B7DE 16'hB74A
`define CUBE_LUT_B7DF 16'hB74B
`define CUBE_LUT_B7E0 16'hB74C
`define CUBE_LUT_B7E1 16'hB74C
`define CUBE_LUT_B7E2 16'hB74D
`define CUBE_LUT_B7E3 16'hB74E
`define CUBE_LUT_B7E4 16'hB74F
`define CUBE_LUT_B7E5 16'hB750
`define CUBE_LUT_B7E6 16'hB750
`define CUBE_LUT_B7E7 16'hB751
`define CUBE_LUT_B7E8 16'hB752
`define CUBE_LUT_B7E9 16'hB753
`define CUBE_LUT_B7EA 16'hB753
`define CUBE_LUT_B7EB 16'hB754
`define CUBE_LUT_B7EC 16'hB755
`define CUBE_LUT_B7ED 16'hB756
`define CUBE_LUT_B7EE 16'hB757
`define CUBE_LUT_B7EF 16'hB757
`define CUBE_LUT_B7F0 16'hB758
`define CUBE_LUT_B7F1 16'hB759
`define CUBE_LUT_B7F2 16'hB75A
`define CUBE_LUT_B7F3 16'hB75B
`define CUBE_LUT_B7F4 16'hB75B
`define CUBE_LUT_B7F5 16'hB75C
`define CUBE_LUT_B7F6 16'hB75D
`define CUBE_LUT_B7F7 16'hB75E
`define CUBE_LUT_B7F8 16'hB75F
`define CUBE_LUT_B7F9 16'hB75F
`define CUBE_LUT_B7FA 16'hB760
`define CUBE_LUT_B7FB 16'hB761
`define CUBE_LUT_B7FC 16'hB762
`define CUBE_LUT_B7FD 16'hB762
`define CUBE_LUT_B7FE 16'hB763
`define CUBE_LUT_B7FF 16'hB764
`define CUBE_LUT_B800 16'hB765
`define CUBE_LUT_B801 16'hB766
`define CUBE_LUT_B802 16'hB768
`define CUBE_LUT_B803 16'hB76A
`define CUBE_LUT_B804 16'hB76B
`define CUBE_LUT_B805 16'hB76D
`define CUBE_LUT_B806 16'hB76E
`define CUBE_LUT_B807 16'hB770
`define CUBE_LUT_B808 16'hB771
`define CUBE_LUT_B809 16'hB773
`define CUBE_LUT_B80A 16'hB775
`define CUBE_LUT_B80B 16'hB776
`define CUBE_LUT_B80C 16'hB778
`define CUBE_LUT_B80D 16'hB779
`define CUBE_LUT_B80E 16'hB77B
`define CUBE_LUT_B80F 16'hB77C
`define CUBE_LUT_B810 16'hB77E
`define CUBE_LUT_B811 16'hB77F
`define CUBE_LUT_B812 16'hB781
`define CUBE_LUT_B813 16'hB783
`define CUBE_LUT_B814 16'hB784
`define CUBE_LUT_B815 16'hB786
`define CUBE_LUT_B816 16'hB787
`define CUBE_LUT_B817 16'hB789
`define CUBE_LUT_B818 16'hB78A
`define CUBE_LUT_B819 16'hB78C
`define CUBE_LUT_B81A 16'hB78D
`define CUBE_LUT_B81B 16'hB78F
`define CUBE_LUT_B81C 16'hB791
`define CUBE_LUT_B81D 16'hB792
`define CUBE_LUT_B81E 16'hB794
`define CUBE_LUT_B81F 16'hB795
`define CUBE_LUT_B820 16'hB797
`define CUBE_LUT_B821 16'hB798
`define CUBE_LUT_B822 16'hB79A
`define CUBE_LUT_B823 16'hB79B
`define CUBE_LUT_B824 16'hB79D
`define CUBE_LUT_B825 16'hB79F
`define CUBE_LUT_B826 16'hB7A0
`define CUBE_LUT_B827 16'hB7A2
`define CUBE_LUT_B828 16'hB7A3
`define CUBE_LUT_B829 16'hB7A5
`define CUBE_LUT_B82A 16'hB7A6
`define CUBE_LUT_B82B 16'hB7A8
`define CUBE_LUT_B82C 16'hB7A9
`define CUBE_LUT_B82D 16'hB7AB
`define CUBE_LUT_B82E 16'hB7AC
`define CUBE_LUT_B82F 16'hB7AE
`define CUBE_LUT_B830 16'hB7B0
`define CUBE_LUT_B831 16'hB7B1
`define CUBE_LUT_B832 16'hB7B3
`define CUBE_LUT_B833 16'hB7B4
`define CUBE_LUT_B834 16'hB7B6
`define CUBE_LUT_B835 16'hB7B7
`define CUBE_LUT_B836 16'hB7B9
`define CUBE_LUT_B837 16'hB7BA
`define CUBE_LUT_B838 16'hB7BC
`define CUBE_LUT_B839 16'hB7BD
`define CUBE_LUT_B83A 16'hB7BF
`define CUBE_LUT_B83B 16'hB7C0
`define CUBE_LUT_B83C 16'hB7C2
`define CUBE_LUT_B83D 16'hB7C3
`define CUBE_LUT_B83E 16'hB7C5
`define CUBE_LUT_B83F 16'hB7C7
`define CUBE_LUT_B840 16'hB7C8
`define CUBE_LUT_B841 16'hB7CA
`define CUBE_LUT_B842 16'hB7CB
`define CUBE_LUT_B843 16'hB7CD
`define CUBE_LUT_B844 16'hB7CE
`define CUBE_LUT_B845 16'hB7D0
`define CUBE_LUT_B846 16'hB7D1
`define CUBE_LUT_B847 16'hB7D3
`define CUBE_LUT_B848 16'hB7D4
`define CUBE_LUT_B849 16'hB7D6
`define CUBE_LUT_B84A 16'hB7D7
`define CUBE_LUT_B84B 16'hB7D9
`define CUBE_LUT_B84C 16'hB7DA
`define CUBE_LUT_B84D 16'hB7DC
`define CUBE_LUT_B84E 16'hB7DD
`define CUBE_LUT_B84F 16'hB7DF
`define CUBE_LUT_B850 16'hB7E0
`define CUBE_LUT_B851 16'hB7E2
`define CUBE_LUT_B852 16'hB7E3
`define CUBE_LUT_B853 16'hB7E5
`define CUBE_LUT_B854 16'hB7E6
`define CUBE_LUT_B855 16'hB7E8
`define CUBE_LUT_B856 16'hB7E9
`define CUBE_LUT_B857 16'hB7EB
`define CUBE_LUT_B858 16'hB7EC
`define CUBE_LUT_B859 16'hB7EE
`define CUBE_LUT_B85A 16'hB7EF
`define CUBE_LUT_B85B 16'hB7F1
`define CUBE_LUT_B85C 16'hB7F3
`define CUBE_LUT_B85D 16'hB7F4
`define CUBE_LUT_B85E 16'hB7F6
`define CUBE_LUT_B85F 16'hB7F7
`define CUBE_LUT_B860 16'hB7F9
`define CUBE_LUT_B861 16'hB7FA
`define CUBE_LUT_B862 16'hB7FC
`define CUBE_LUT_B863 16'hB7FD
`define CUBE_LUT_B864 16'hB7FF
`define CUBE_LUT_B865 16'hB800
`define CUBE_LUT_B866 16'hB801
`define CUBE_LUT_B867 16'hB802
`define CUBE_LUT_B868 16'hB802
`define CUBE_LUT_B869 16'hB803
`define CUBE_LUT_B86A 16'hB804
`define CUBE_LUT_B86B 16'hB805
`define CUBE_LUT_B86C 16'hB805
`define CUBE_LUT_B86D 16'hB806
`define CUBE_LUT_B86E 16'hB807
`define CUBE_LUT_B86F 16'hB807
`define CUBE_LUT_B870 16'hB808
`define CUBE_LUT_B871 16'hB809
`define CUBE_LUT_B872 16'hB80A
`define CUBE_LUT_B873 16'hB80A
`define CUBE_LUT_B874 16'hB80B
`define CUBE_LUT_B875 16'hB80C
`define CUBE_LUT_B876 16'hB80D
`define CUBE_LUT_B877 16'hB80D
`define CUBE_LUT_B878 16'hB80E
`define CUBE_LUT_B879 16'hB80F
`define CUBE_LUT_B87A 16'hB810
`define CUBE_LUT_B87B 16'hB810
`define CUBE_LUT_B87C 16'hB811
`define CUBE_LUT_B87D 16'hB812
`define CUBE_LUT_B87E 16'hB813
`define CUBE_LUT_B87F 16'hB813
`define CUBE_LUT_B880 16'hB814
`define CUBE_LUT_B881 16'hB815
`define CUBE_LUT_B882 16'hB816
`define CUBE_LUT_B883 16'hB816
`define CUBE_LUT_B884 16'hB817
`define CUBE_LUT_B885 16'hB818
`define CUBE_LUT_B886 16'hB819
`define CUBE_LUT_B887 16'hB819
`define CUBE_LUT_B888 16'hB81A
`define CUBE_LUT_B889 16'hB81B
`define CUBE_LUT_B88A 16'hB81C
`define CUBE_LUT_B88B 16'hB81C
`define CUBE_LUT_B88C 16'hB81D
`define CUBE_LUT_B88D 16'hB81E
`define CUBE_LUT_B88E 16'hB81E
`define CUBE_LUT_B88F 16'hB81F
`define CUBE_LUT_B890 16'hB820
`define CUBE_LUT_B891 16'hB821
`define CUBE_LUT_B892 16'hB821
`define CUBE_LUT_B893 16'hB822
`define CUBE_LUT_B894 16'hB823
`define CUBE_LUT_B895 16'hB824
`define CUBE_LUT_B896 16'hB824
`define CUBE_LUT_B897 16'hB825
`define CUBE_LUT_B898 16'hB826
`define CUBE_LUT_B899 16'hB827
`define CUBE_LUT_B89A 16'hB827
`define CUBE_LUT_B89B 16'hB828
`define CUBE_LUT_B89C 16'hB829
`define CUBE_LUT_B89D 16'hB829
`define CUBE_LUT_B89E 16'hB82A
`define CUBE_LUT_B89F 16'hB82B
`define CUBE_LUT_B8A0 16'hB82C
`define CUBE_LUT_B8A1 16'hB82C
`define CUBE_LUT_B8A2 16'hB82D
`define CUBE_LUT_B8A3 16'hB82E
`define CUBE_LUT_B8A4 16'hB82F
`define CUBE_LUT_B8A5 16'hB82F
`define CUBE_LUT_B8A6 16'hB830
`define CUBE_LUT_B8A7 16'hB831
`define CUBE_LUT_B8A8 16'hB831
`define CUBE_LUT_B8A9 16'hB832
`define CUBE_LUT_B8AA 16'hB833
`define CUBE_LUT_B8AB 16'hB834
`define CUBE_LUT_B8AC 16'hB834
`define CUBE_LUT_B8AD 16'hB835
`define CUBE_LUT_B8AE 16'hB836
`define CUBE_LUT_B8AF 16'hB837
`define CUBE_LUT_B8B0 16'hB837
`define CUBE_LUT_B8B1 16'hB838
`define CUBE_LUT_B8B2 16'hB839
`define CUBE_LUT_B8B3 16'hB839
`define CUBE_LUT_B8B4 16'hB83A
`define CUBE_LUT_B8B5 16'hB83B
`define CUBE_LUT_B8B6 16'hB83C
`define CUBE_LUT_B8B7 16'hB83C
`define CUBE_LUT_B8B8 16'hB83D
`define CUBE_LUT_B8B9 16'hB83E
`define CUBE_LUT_B8BA 16'hB83E
`define CUBE_LUT_B8BB 16'hB83F
`define CUBE_LUT_B8BC 16'hB840
`define CUBE_LUT_B8BD 16'hB841
`define CUBE_LUT_B8BE 16'hB841
`define CUBE_LUT_B8BF 16'hB842
`define CUBE_LUT_B8C0 16'hB843
`define CUBE_LUT_B8C1 16'hB843
`define CUBE_LUT_B8C2 16'hB844
`define CUBE_LUT_B8C3 16'hB845
`define CUBE_LUT_B8C4 16'hB846
`define CUBE_LUT_B8C5 16'hB846
`define CUBE_LUT_B8C6 16'hB847
`define CUBE_LUT_B8C7 16'hB848
`define CUBE_LUT_B8C8 16'hB848
`define CUBE_LUT_B8C9 16'hB849
`define CUBE_LUT_B8CA 16'hB84A
`define CUBE_LUT_B8CB 16'hB84B
`define CUBE_LUT_B8CC 16'hB84B
`define CUBE_LUT_B8CD 16'hB84C
`define CUBE_LUT_B8CE 16'hB84D
`define CUBE_LUT_B8CF 16'hB84D
`define CUBE_LUT_B8D0 16'hB84E
`define CUBE_LUT_B8D1 16'hB84F
`define CUBE_LUT_B8D2 16'hB850
`define CUBE_LUT_B8D3 16'hB850
`define CUBE_LUT_B8D4 16'hB851
`define CUBE_LUT_B8D5 16'hB852
`define CUBE_LUT_B8D6 16'hB852
`define CUBE_LUT_B8D7 16'hB853
`define CUBE_LUT_B8D8 16'hB854
`define CUBE_LUT_B8D9 16'hB855
`define CUBE_LUT_B8DA 16'hB855
`define CUBE_LUT_B8DB 16'hB856
`define CUBE_LUT_B8DC 16'hB857
`define CUBE_LUT_B8DD 16'hB857
`define CUBE_LUT_B8DE 16'hB858
`define CUBE_LUT_B8DF 16'hB859
`define CUBE_LUT_B8E0 16'hB859
`define CUBE_LUT_B8E1 16'hB85A
`define CUBE_LUT_B8E2 16'hB85B
`define CUBE_LUT_B8E3 16'hB85C
`define CUBE_LUT_B8E4 16'hB85C
`define CUBE_LUT_B8E5 16'hB85D
`define CUBE_LUT_B8E6 16'hB85E
`define CUBE_LUT_B8E7 16'hB85E
`define CUBE_LUT_B8E8 16'hB85F
`define CUBE_LUT_B8E9 16'hB860
`define CUBE_LUT_B8EA 16'hB860
`define CUBE_LUT_B8EB 16'hB861
`define CUBE_LUT_B8EC 16'hB862
`define CUBE_LUT_B8ED 16'hB863
`define CUBE_LUT_B8EE 16'hB863
`define CUBE_LUT_B8EF 16'hB864
`define CUBE_LUT_B8F0 16'hB865
`define CUBE_LUT_B8F1 16'hB865
`define CUBE_LUT_B8F2 16'hB866
`define CUBE_LUT_B8F3 16'hB867
`define CUBE_LUT_B8F4 16'hB867
`define CUBE_LUT_B8F5 16'hB868
`define CUBE_LUT_B8F6 16'hB869
`define CUBE_LUT_B8F7 16'hB86A
`define CUBE_LUT_B8F8 16'hB86A
`define CUBE_LUT_B8F9 16'hB86B
`define CUBE_LUT_B8FA 16'hB86C
`define CUBE_LUT_B8FB 16'hB86C
`define CUBE_LUT_B8FC 16'hB86D
`define CUBE_LUT_B8FD 16'hB86E
`define CUBE_LUT_B8FE 16'hB86E
`define CUBE_LUT_B8FF 16'hB86F
`define CUBE_LUT_B900 16'hB870
`define CUBE_LUT_B901 16'hB871
`define CUBE_LUT_B902 16'hB871
`define CUBE_LUT_B903 16'hB872
`define CUBE_LUT_B904 16'hB873
`define CUBE_LUT_B905 16'hB873
`define CUBE_LUT_B906 16'hB874
`define CUBE_LUT_B907 16'hB875
`define CUBE_LUT_B908 16'hB875
`define CUBE_LUT_B909 16'hB876
`define CUBE_LUT_B90A 16'hB877
`define CUBE_LUT_B90B 16'hB877
`define CUBE_LUT_B90C 16'hB878
`define CUBE_LUT_B90D 16'hB879
`define CUBE_LUT_B90E 16'hB879
`define CUBE_LUT_B90F 16'hB87A
`define CUBE_LUT_B910 16'hB87B
`define CUBE_LUT_B911 16'hB87C
`define CUBE_LUT_B912 16'hB87C
`define CUBE_LUT_B913 16'hB87D
`define CUBE_LUT_B914 16'hB87E
`define CUBE_LUT_B915 16'hB87E
`define CUBE_LUT_B916 16'hB87F
`define CUBE_LUT_B917 16'hB880
`define CUBE_LUT_B918 16'hB880
`define CUBE_LUT_B919 16'hB881
`define CUBE_LUT_B91A 16'hB882
`define CUBE_LUT_B91B 16'hB882
`define CUBE_LUT_B91C 16'hB883
`define CUBE_LUT_B91D 16'hB884
`define CUBE_LUT_B91E 16'hB884
`define CUBE_LUT_B91F 16'hB885
`define CUBE_LUT_B920 16'hB886
`define CUBE_LUT_B921 16'hB886
`define CUBE_LUT_B922 16'hB887
`define CUBE_LUT_B923 16'hB888
`define CUBE_LUT_B924 16'hB889
`define CUBE_LUT_B925 16'hB889
`define CUBE_LUT_B926 16'hB88A
`define CUBE_LUT_B927 16'hB88B
`define CUBE_LUT_B928 16'hB88B
`define CUBE_LUT_B929 16'hB88C
`define CUBE_LUT_B92A 16'hB88D
`define CUBE_LUT_B92B 16'hB88D
`define CUBE_LUT_B92C 16'hB88E
`define CUBE_LUT_B92D 16'hB88F
`define CUBE_LUT_B92E 16'hB88F
`define CUBE_LUT_B92F 16'hB890
`define CUBE_LUT_B930 16'hB891
`define CUBE_LUT_B931 16'hB891
`define CUBE_LUT_B932 16'hB892
`define CUBE_LUT_B933 16'hB893
`define CUBE_LUT_B934 16'hB893
`define CUBE_LUT_B935 16'hB894
`define CUBE_LUT_B936 16'hB895
`define CUBE_LUT_B937 16'hB895
`define CUBE_LUT_B938 16'hB896
`define CUBE_LUT_B939 16'hB897
`define CUBE_LUT_B93A 16'hB897
`define CUBE_LUT_B93B 16'hB898
`define CUBE_LUT_B93C 16'hB899
`define CUBE_LUT_B93D 16'hB899
`define CUBE_LUT_B93E 16'hB89A
`define CUBE_LUT_B93F 16'hB89B
`define CUBE_LUT_B940 16'hB89B
`define CUBE_LUT_B941 16'hB89C
`define CUBE_LUT_B942 16'hB89D
`define CUBE_LUT_B943 16'hB89D
`define CUBE_LUT_B944 16'hB89E
`define CUBE_LUT_B945 16'hB89F
`define CUBE_LUT_B946 16'hB89F
`define CUBE_LUT_B947 16'hB8A0
`define CUBE_LUT_B948 16'hB8A1
`define CUBE_LUT_B949 16'hB8A1
`define CUBE_LUT_B94A 16'hB8A2
`define CUBE_LUT_B94B 16'hB8A3
`define CUBE_LUT_B94C 16'hB8A3
`define CUBE_LUT_B94D 16'hB8A4
`define CUBE_LUT_B94E 16'hB8A5
`define CUBE_LUT_B94F 16'hB8A5
`define CUBE_LUT_B950 16'hB8A6
`define CUBE_LUT_B951 16'hB8A7
`define CUBE_LUT_B952 16'hB8A7
`define CUBE_LUT_B953 16'hB8A8
`define CUBE_LUT_B954 16'hB8A9
`define CUBE_LUT_B955 16'hB8A9
`define CUBE_LUT_B956 16'hB8AA
`define CUBE_LUT_B957 16'hB8AB
`define CUBE_LUT_B958 16'hB8AB
`define CUBE_LUT_B959 16'hB8AC
`define CUBE_LUT_B95A 16'hB8AD
`define CUBE_LUT_B95B 16'hB8AD
`define CUBE_LUT_B95C 16'hB8AE
`define CUBE_LUT_B95D 16'hB8AF
`define CUBE_LUT_B95E 16'hB8AF
`define CUBE_LUT_B95F 16'hB8B0
`define CUBE_LUT_B960 16'hB8B1
`define CUBE_LUT_B961 16'hB8B1
`define CUBE_LUT_B962 16'hB8B2
`define CUBE_LUT_B963 16'hB8B3
`define CUBE_LUT_B964 16'hB8B3
`define CUBE_LUT_B965 16'hB8B4
`define CUBE_LUT_B966 16'hB8B4
`define CUBE_LUT_B967 16'hB8B5
`define CUBE_LUT_B968 16'hB8B6
`define CUBE_LUT_B969 16'hB8B6
`define CUBE_LUT_B96A 16'hB8B7
`define CUBE_LUT_B96B 16'hB8B8
`define CUBE_LUT_B96C 16'hB8B8
`define CUBE_LUT_B96D 16'hB8B9
`define CUBE_LUT_B96E 16'hB8BA
`define CUBE_LUT_B96F 16'hB8BA
`define CUBE_LUT_B970 16'hB8BB
`define CUBE_LUT_B971 16'hB8BC
`define CUBE_LUT_B972 16'hB8BC
`define CUBE_LUT_B973 16'hB8BD
`define CUBE_LUT_B974 16'hB8BE
`define CUBE_LUT_B975 16'hB8BE
`define CUBE_LUT_B976 16'hB8BF
`define CUBE_LUT_B977 16'hB8C0
`define CUBE_LUT_B978 16'hB8C0
`define CUBE_LUT_B979 16'hB8C1
`define CUBE_LUT_B97A 16'hB8C2
`define CUBE_LUT_B97B 16'hB8C2
`define CUBE_LUT_B97C 16'hB8C3
`define CUBE_LUT_B97D 16'hB8C3
`define CUBE_LUT_B97E 16'hB8C4
`define CUBE_LUT_B97F 16'hB8C5
`define CUBE_LUT_B980 16'hB8C5
`define CUBE_LUT_B981 16'hB8C6
`define CUBE_LUT_B982 16'hB8C7
`define CUBE_LUT_B983 16'hB8C7
`define CUBE_LUT_B984 16'hB8C8
`define CUBE_LUT_B985 16'hB8C9
`define CUBE_LUT_B986 16'hB8C9
`define CUBE_LUT_B987 16'hB8CA
`define CUBE_LUT_B988 16'hB8CB
`define CUBE_LUT_B989 16'hB8CB
`define CUBE_LUT_B98A 16'hB8CC
`define CUBE_LUT_B98B 16'hB8CC
`define CUBE_LUT_B98C 16'hB8CD
`define CUBE_LUT_B98D 16'hB8CE
`define CUBE_LUT_B98E 16'hB8CE
`define CUBE_LUT_B98F 16'hB8CF
`define CUBE_LUT_B990 16'hB8D0
`define CUBE_LUT_B991 16'hB8D0
`define CUBE_LUT_B992 16'hB8D1
`define CUBE_LUT_B993 16'hB8D2
`define CUBE_LUT_B994 16'hB8D2
`define CUBE_LUT_B995 16'hB8D3
`define CUBE_LUT_B996 16'hB8D3
`define CUBE_LUT_B997 16'hB8D4
`define CUBE_LUT_B998 16'hB8D5
`define CUBE_LUT_B999 16'hB8D5
`define CUBE_LUT_B99A 16'hB8D6
`define CUBE_LUT_B99B 16'hB8D7
`define CUBE_LUT_B99C 16'hB8D7
`define CUBE_LUT_B99D 16'hB8D8
`define CUBE_LUT_B99E 16'hB8D9
`define CUBE_LUT_B99F 16'hB8D9
`define CUBE_LUT_B9A0 16'hB8DA
`define CUBE_LUT_B9A1 16'hB8DA
`define CUBE_LUT_B9A2 16'hB8DB
`define CUBE_LUT_B9A3 16'hB8DC
`define CUBE_LUT_B9A4 16'hB8DC
`define CUBE_LUT_B9A5 16'hB8DD
`define CUBE_LUT_B9A6 16'hB8DE
`define CUBE_LUT_B9A7 16'hB8DE
`define CUBE_LUT_B9A8 16'hB8DF
`define CUBE_LUT_B9A9 16'hB8DF
`define CUBE_LUT_B9AA 16'hB8E0
`define CUBE_LUT_B9AB 16'hB8E1
`define CUBE_LUT_B9AC 16'hB8E1
`define CUBE_LUT_B9AD 16'hB8E2
`define CUBE_LUT_B9AE 16'hB8E3
`define CUBE_LUT_B9AF 16'hB8E3
`define CUBE_LUT_B9B0 16'hB8E4
`define CUBE_LUT_B9B1 16'hB8E4
`define CUBE_LUT_B9B2 16'hB8E5
`define CUBE_LUT_B9B3 16'hB8E6
`define CUBE_LUT_B9B4 16'hB8E6
`define CUBE_LUT_B9B5 16'hB8E7
`define CUBE_LUT_B9B6 16'hB8E8
`define CUBE_LUT_B9B7 16'hB8E8
`define CUBE_LUT_B9B8 16'hB8E9
`define CUBE_LUT_B9B9 16'hB8E9
`define CUBE_LUT_B9BA 16'hB8EA
`define CUBE_LUT_B9BB 16'hB8EB
`define CUBE_LUT_B9BC 16'hB8EB
`define CUBE_LUT_B9BD 16'hB8EC
`define CUBE_LUT_B9BE 16'hB8ED
`define CUBE_LUT_B9BF 16'hB8ED
`define CUBE_LUT_B9C0 16'hB8EE
`define CUBE_LUT_B9C1 16'hB8EE
`define CUBE_LUT_B9C2 16'hB8EF
`define CUBE_LUT_B9C3 16'hB8F0
`define CUBE_LUT_B9C4 16'hB8F0
`define CUBE_LUT_B9C5 16'hB8F1
`define CUBE_LUT_B9C6 16'hB8F2
`define CUBE_LUT_B9C7 16'hB8F2
`define CUBE_LUT_B9C8 16'hB8F3
`define CUBE_LUT_B9C9 16'hB8F3
`define CUBE_LUT_B9CA 16'hB8F4
`define CUBE_LUT_B9CB 16'hB8F5
`define CUBE_LUT_B9CC 16'hB8F5
`define CUBE_LUT_B9CD 16'hB8F6
`define CUBE_LUT_B9CE 16'hB8F6
`define CUBE_LUT_B9CF 16'hB8F7
`define CUBE_LUT_B9D0 16'hB8F8
`define CUBE_LUT_B9D1 16'hB8F8
`define CUBE_LUT_B9D2 16'hB8F9
`define CUBE_LUT_B9D3 16'hB8FA
`define CUBE_LUT_B9D4 16'hB8FA
`define CUBE_LUT_B9D5 16'hB8FB
`define CUBE_LUT_B9D6 16'hB8FB
`define CUBE_LUT_B9D7 16'hB8FC
`define CUBE_LUT_B9D8 16'hB8FD
`define CUBE_LUT_B9D9 16'hB8FD
`define CUBE_LUT_B9DA 16'hB8FE
`define CUBE_LUT_B9DB 16'hB8FE
`define CUBE_LUT_B9DC 16'hB8FF
`define CUBE_LUT_B9DD 16'hB900
`define CUBE_LUT_B9DE 16'hB900
`define CUBE_LUT_B9DF 16'hB901
`define CUBE_LUT_B9E0 16'hB902
`define CUBE_LUT_B9E1 16'hB902
`define CUBE_LUT_B9E2 16'hB903
`define CUBE_LUT_B9E3 16'hB903
`define CUBE_LUT_B9E4 16'hB904
`define CUBE_LUT_B9E5 16'hB905
`define CUBE_LUT_B9E6 16'hB905
`define CUBE_LUT_B9E7 16'hB906
`define CUBE_LUT_B9E8 16'hB906
`define CUBE_LUT_B9E9 16'hB907
`define CUBE_LUT_B9EA 16'hB908
`define CUBE_LUT_B9EB 16'hB908
`define CUBE_LUT_B9EC 16'hB909
`define CUBE_LUT_B9ED 16'hB909
`define CUBE_LUT_B9EE 16'hB90A
`define CUBE_LUT_B9EF 16'hB90B
`define CUBE_LUT_B9F0 16'hB90B
`define CUBE_LUT_B9F1 16'hB90C
`define CUBE_LUT_B9F2 16'hB90C
`define CUBE_LUT_B9F3 16'hB90D
`define CUBE_LUT_B9F4 16'hB90E
`define CUBE_LUT_B9F5 16'hB90E
`define CUBE_LUT_B9F6 16'hB90F
`define CUBE_LUT_B9F7 16'hB90F
`define CUBE_LUT_B9F8 16'hB910
`define CUBE_LUT_B9F9 16'hB911
`define CUBE_LUT_B9FA 16'hB911
`define CUBE_LUT_B9FB 16'hB912
`define CUBE_LUT_B9FC 16'hB912
`define CUBE_LUT_B9FD 16'hB913
`define CUBE_LUT_B9FE 16'hB914
`define CUBE_LUT_B9FF 16'hB914
`define CUBE_LUT_BA00 16'hB915
`define CUBE_LUT_BA01 16'hB915
`define CUBE_LUT_BA02 16'hB916
`define CUBE_LUT_BA03 16'hB917
`define CUBE_LUT_BA04 16'hB917
`define CUBE_LUT_BA05 16'hB918
`define CUBE_LUT_BA06 16'hB918
`define CUBE_LUT_BA07 16'hB919
`define CUBE_LUT_BA08 16'hB91A
`define CUBE_LUT_BA09 16'hB91A
`define CUBE_LUT_BA0A 16'hB91B
`define CUBE_LUT_BA0B 16'hB91B
`define CUBE_LUT_BA0C 16'hB91C
`define CUBE_LUT_BA0D 16'hB91D
`define CUBE_LUT_BA0E 16'hB91D
`define CUBE_LUT_BA0F 16'hB91E
`define CUBE_LUT_BA10 16'hB91E
`define CUBE_LUT_BA11 16'hB91F
`define CUBE_LUT_BA12 16'hB91F
`define CUBE_LUT_BA13 16'hB920
`define CUBE_LUT_BA14 16'hB921
`define CUBE_LUT_BA15 16'hB921
`define CUBE_LUT_BA16 16'hB922
`define CUBE_LUT_BA17 16'hB922
`define CUBE_LUT_BA18 16'hB923
`define CUBE_LUT_BA19 16'hB924
`define CUBE_LUT_BA1A 16'hB924
`define CUBE_LUT_BA1B 16'hB925
`define CUBE_LUT_BA1C 16'hB925
`define CUBE_LUT_BA1D 16'hB926
`define CUBE_LUT_BA1E 16'hB927
`define CUBE_LUT_BA1F 16'hB927
`define CUBE_LUT_BA20 16'hB928
`define CUBE_LUT_BA21 16'hB928
`define CUBE_LUT_BA22 16'hB929
`define CUBE_LUT_BA23 16'hB929
`define CUBE_LUT_BA24 16'hB92A
`define CUBE_LUT_BA25 16'hB92B
`define CUBE_LUT_BA26 16'hB92B
`define CUBE_LUT_BA27 16'hB92C
`define CUBE_LUT_BA28 16'hB92C
`define CUBE_LUT_BA29 16'hB92D
`define CUBE_LUT_BA2A 16'hB92E
`define CUBE_LUT_BA2B 16'hB92E
`define CUBE_LUT_BA2C 16'hB92F
`define CUBE_LUT_BA2D 16'hB92F
`define CUBE_LUT_BA2E 16'hB930
`define CUBE_LUT_BA2F 16'hB930
`define CUBE_LUT_BA30 16'hB931
`define CUBE_LUT_BA31 16'hB932
`define CUBE_LUT_BA32 16'hB932
`define CUBE_LUT_BA33 16'hB933
`define CUBE_LUT_BA34 16'hB933
`define CUBE_LUT_BA35 16'hB934
`define CUBE_LUT_BA36 16'hB934
`define CUBE_LUT_BA37 16'hB935
`define CUBE_LUT_BA38 16'hB936
`define CUBE_LUT_BA39 16'hB936
`define CUBE_LUT_BA3A 16'hB937
`define CUBE_LUT_BA3B 16'hB937
`define CUBE_LUT_BA3C 16'hB938
`define CUBE_LUT_BA3D 16'hB938
`define CUBE_LUT_BA3E 16'hB939
`define CUBE_LUT_BA3F 16'hB93A
`define CUBE_LUT_BA40 16'hB93A
`define CUBE_LUT_BA41 16'hB93B
`define CUBE_LUT_BA42 16'hB93B
`define CUBE_LUT_BA43 16'hB93C
`define CUBE_LUT_BA44 16'hB93D
`define CUBE_LUT_BA45 16'hB93D
`define CUBE_LUT_BA46 16'hB93E
`define CUBE_LUT_BA47 16'hB93E
`define CUBE_LUT_BA48 16'hB93F
`define CUBE_LUT_BA49 16'hB93F
`define CUBE_LUT_BA4A 16'hB940
`define CUBE_LUT_BA4B 16'hB940
`define CUBE_LUT_BA4C 16'hB941
`define CUBE_LUT_BA4D 16'hB942
`define CUBE_LUT_BA4E 16'hB942
`define CUBE_LUT_BA4F 16'hB943
`define CUBE_LUT_BA50 16'hB943
`define CUBE_LUT_BA51 16'hB944
`define CUBE_LUT_BA52 16'hB944
`define CUBE_LUT_BA53 16'hB945
`define CUBE_LUT_BA54 16'hB946
`define CUBE_LUT_BA55 16'hB946
`define CUBE_LUT_BA56 16'hB947
`define CUBE_LUT_BA57 16'hB947
`define CUBE_LUT_BA58 16'hB948
`define CUBE_LUT_BA59 16'hB948
`define CUBE_LUT_BA5A 16'hB949
`define CUBE_LUT_BA5B 16'hB94A
`define CUBE_LUT_BA5C 16'hB94A
`define CUBE_LUT_BA5D 16'hB94B
`define CUBE_LUT_BA5E 16'hB94B
`define CUBE_LUT_BA5F 16'hB94C
`define CUBE_LUT_BA60 16'hB94C
`define CUBE_LUT_BA61 16'hB94D
`define CUBE_LUT_BA62 16'hB94D
`define CUBE_LUT_BA63 16'hB94E
`define CUBE_LUT_BA64 16'hB94F
`define CUBE_LUT_BA65 16'hB94F
`define CUBE_LUT_BA66 16'hB950
`define CUBE_LUT_BA67 16'hB950
`define CUBE_LUT_BA68 16'hB951
`define CUBE_LUT_BA69 16'hB951
`define CUBE_LUT_BA6A 16'hB952
`define CUBE_LUT_BA6B 16'hB953
`define CUBE_LUT_BA6C 16'hB953
`define CUBE_LUT_BA6D 16'hB954
`define CUBE_LUT_BA6E 16'hB954
`define CUBE_LUT_BA6F 16'hB955
`define CUBE_LUT_BA70 16'hB955
`define CUBE_LUT_BA71 16'hB956
`define CUBE_LUT_BA72 16'hB956
`define CUBE_LUT_BA73 16'hB957
`define CUBE_LUT_BA74 16'hB958
`define CUBE_LUT_BA75 16'hB958
`define CUBE_LUT_BA76 16'hB959
`define CUBE_LUT_BA77 16'hB959
`define CUBE_LUT_BA78 16'hB95A
`define CUBE_LUT_BA79 16'hB95A
`define CUBE_LUT_BA7A 16'hB95B
`define CUBE_LUT_BA7B 16'hB95B
`define CUBE_LUT_BA7C 16'hB95C
`define CUBE_LUT_BA7D 16'hB95C
`define CUBE_LUT_BA7E 16'hB95D
`define CUBE_LUT_BA7F 16'hB95E
`define CUBE_LUT_BA80 16'hB95E
`define CUBE_LUT_BA81 16'hB95F
`define CUBE_LUT_BA82 16'hB95F
`define CUBE_LUT_BA83 16'hB960
`define CUBE_LUT_BA84 16'hB960
`define CUBE_LUT_BA85 16'hB961
`define CUBE_LUT_BA86 16'hB961
`define CUBE_LUT_BA87 16'hB962
`define CUBE_LUT_BA88 16'hB963
`define CUBE_LUT_BA89 16'hB963
`define CUBE_LUT_BA8A 16'hB964
`define CUBE_LUT_BA8B 16'hB964
`define CUBE_LUT_BA8C 16'hB965
`define CUBE_LUT_BA8D 16'hB965
`define CUBE_LUT_BA8E 16'hB966
`define CUBE_LUT_BA8F 16'hB966
`define CUBE_LUT_BA90 16'hB967
`define CUBE_LUT_BA91 16'hB967
`define CUBE_LUT_BA92 16'hB968
`define CUBE_LUT_BA93 16'hB969
`define CUBE_LUT_BA94 16'hB969
`define CUBE_LUT_BA95 16'hB96A
`define CUBE_LUT_BA96 16'hB96A
`define CUBE_LUT_BA97 16'hB96B
`define CUBE_LUT_BA98 16'hB96B
`define CUBE_LUT_BA99 16'hB96C
`define CUBE_LUT_BA9A 16'hB96C
`define CUBE_LUT_BA9B 16'hB96D
`define CUBE_LUT_BA9C 16'hB96D
`define CUBE_LUT_BA9D 16'hB96E
`define CUBE_LUT_BA9E 16'hB96E
`define CUBE_LUT_BA9F 16'hB96F
`define CUBE_LUT_BAA0 16'hB970
`define CUBE_LUT_BAA1 16'hB970
`define CUBE_LUT_BAA2 16'hB971
`define CUBE_LUT_BAA3 16'hB971
`define CUBE_LUT_BAA4 16'hB972
`define CUBE_LUT_BAA5 16'hB972
`define CUBE_LUT_BAA6 16'hB973
`define CUBE_LUT_BAA7 16'hB973
`define CUBE_LUT_BAA8 16'hB974
`define CUBE_LUT_BAA9 16'hB974
`define CUBE_LUT_BAAA 16'hB975
`define CUBE_LUT_BAAB 16'hB975
`define CUBE_LUT_BAAC 16'hB976
`define CUBE_LUT_BAAD 16'hB977
`define CUBE_LUT_BAAE 16'hB977
`define CUBE_LUT_BAAF 16'hB978
`define CUBE_LUT_BAB0 16'hB978
`define CUBE_LUT_BAB1 16'hB979
`define CUBE_LUT_BAB2 16'hB979
`define CUBE_LUT_BAB3 16'hB97A
`define CUBE_LUT_BAB4 16'hB97A
`define CUBE_LUT_BAB5 16'hB97B
`define CUBE_LUT_BAB6 16'hB97B
`define CUBE_LUT_BAB7 16'hB97C
`define CUBE_LUT_BAB8 16'hB97C
`define CUBE_LUT_BAB9 16'hB97D
`define CUBE_LUT_BABA 16'hB97D
`define CUBE_LUT_BABB 16'hB97E
`define CUBE_LUT_BABC 16'hB97E
`define CUBE_LUT_BABD 16'hB97F
`define CUBE_LUT_BABE 16'hB980
`define CUBE_LUT_BABF 16'hB980
`define CUBE_LUT_BAC0 16'hB981
`define CUBE_LUT_BAC1 16'hB981
`define CUBE_LUT_BAC2 16'hB982
`define CUBE_LUT_BAC3 16'hB982
`define CUBE_LUT_BAC4 16'hB983
`define CUBE_LUT_BAC5 16'hB983
`define CUBE_LUT_BAC6 16'hB984
`define CUBE_LUT_BAC7 16'hB984
`define CUBE_LUT_BAC8 16'hB985
`define CUBE_LUT_BAC9 16'hB985
`define CUBE_LUT_BACA 16'hB986
`define CUBE_LUT_BACB 16'hB986
`define CUBE_LUT_BACC 16'hB987
`define CUBE_LUT_BACD 16'hB987
`define CUBE_LUT_BACE 16'hB988
`define CUBE_LUT_BACF 16'hB988
`define CUBE_LUT_BAD0 16'hB989
`define CUBE_LUT_BAD1 16'hB98A
`define CUBE_LUT_BAD2 16'hB98A
`define CUBE_LUT_BAD3 16'hB98B
`define CUBE_LUT_BAD4 16'hB98B
`define CUBE_LUT_BAD5 16'hB98C
`define CUBE_LUT_BAD6 16'hB98C
`define CUBE_LUT_BAD7 16'hB98D
`define CUBE_LUT_BAD8 16'hB98D
`define CUBE_LUT_BAD9 16'hB98E
`define CUBE_LUT_BADA 16'hB98E
`define CUBE_LUT_BADB 16'hB98F
`define CUBE_LUT_BADC 16'hB98F
`define CUBE_LUT_BADD 16'hB990
`define CUBE_LUT_BADE 16'hB990
`define CUBE_LUT_BADF 16'hB991
`define CUBE_LUT_BAE0 16'hB991
`define CUBE_LUT_BAE1 16'hB992
`define CUBE_LUT_BAE2 16'hB992
`define CUBE_LUT_BAE3 16'hB993
`define CUBE_LUT_BAE4 16'hB993
`define CUBE_LUT_BAE5 16'hB994
`define CUBE_LUT_BAE6 16'hB994
`define CUBE_LUT_BAE7 16'hB995
`define CUBE_LUT_BAE8 16'hB995
`define CUBE_LUT_BAE9 16'hB996
`define CUBE_LUT_BAEA 16'hB996
`define CUBE_LUT_BAEB 16'hB997
`define CUBE_LUT_BAEC 16'hB997
`define CUBE_LUT_BAED 16'hB998
`define CUBE_LUT_BAEE 16'hB998
`define CUBE_LUT_BAEF 16'hB999
`define CUBE_LUT_BAF0 16'hB999
`define CUBE_LUT_BAF1 16'hB99A
`define CUBE_LUT_BAF2 16'hB99B
`define CUBE_LUT_BAF3 16'hB99B
`define CUBE_LUT_BAF4 16'hB99C
`define CUBE_LUT_BAF5 16'hB99C
`define CUBE_LUT_BAF6 16'hB99D
`define CUBE_LUT_BAF7 16'hB99D
`define CUBE_LUT_BAF8 16'hB99E
`define CUBE_LUT_BAF9 16'hB99E
`define CUBE_LUT_BAFA 16'hB99F
`define CUBE_LUT_BAFB 16'hB99F
`define CUBE_LUT_BAFC 16'hB9A0
`define CUBE_LUT_BAFD 16'hB9A0
`define CUBE_LUT_BAFE 16'hB9A1
`define CUBE_LUT_BAFF 16'hB9A1
`define CUBE_LUT_BB00 16'hB9A2
`define CUBE_LUT_BB01 16'hB9A2
`define CUBE_LUT_BB02 16'hB9A3
`define CUBE_LUT_BB03 16'hB9A3
`define CUBE_LUT_BB04 16'hB9A4
`define CUBE_LUT_BB05 16'hB9A4
`define CUBE_LUT_BB06 16'hB9A5
`define CUBE_LUT_BB07 16'hB9A5
`define CUBE_LUT_BB08 16'hB9A6
`define CUBE_LUT_BB09 16'hB9A6
`define CUBE_LUT_BB0A 16'hB9A7
`define CUBE_LUT_BB0B 16'hB9A7
`define CUBE_LUT_BB0C 16'hB9A8
`define CUBE_LUT_BB0D 16'hB9A8
`define CUBE_LUT_BB0E 16'hB9A9
`define CUBE_LUT_BB0F 16'hB9A9
`define CUBE_LUT_BB10 16'hB9AA
`define CUBE_LUT_BB11 16'hB9AA
`define CUBE_LUT_BB12 16'hB9AB
`define CUBE_LUT_BB13 16'hB9AB
`define CUBE_LUT_BB14 16'hB9AC
`define CUBE_LUT_BB15 16'hB9AC
`define CUBE_LUT_BB16 16'hB9AD
`define CUBE_LUT_BB17 16'hB9AD
`define CUBE_LUT_BB18 16'hB9AE
`define CUBE_LUT_BB19 16'hB9AE
`define CUBE_LUT_BB1A 16'hB9AF
`define CUBE_LUT_BB1B 16'hB9AF
`define CUBE_LUT_BB1C 16'hB9B0
`define CUBE_LUT_BB1D 16'hB9B0
`define CUBE_LUT_BB1E 16'hB9B1
`define CUBE_LUT_BB1F 16'hB9B1
`define CUBE_LUT_BB20 16'hB9B2
`define CUBE_LUT_BB21 16'hB9B2
`define CUBE_LUT_BB22 16'hB9B3
`define CUBE_LUT_BB23 16'hB9B3
`define CUBE_LUT_BB24 16'hB9B4
`define CUBE_LUT_BB25 16'hB9B4
`define CUBE_LUT_BB26 16'hB9B5
`define CUBE_LUT_BB27 16'hB9B5
`define CUBE_LUT_BB28 16'hB9B6
`define CUBE_LUT_BB29 16'hB9B6
`define CUBE_LUT_BB2A 16'hB9B6
`define CUBE_LUT_BB2B 16'hB9B7
`define CUBE_LUT_BB2C 16'hB9B7
`define CUBE_LUT_BB2D 16'hB9B8
`define CUBE_LUT_BB2E 16'hB9B8
`define CUBE_LUT_BB2F 16'hB9B9
`define CUBE_LUT_BB30 16'hB9B9
`define CUBE_LUT_BB31 16'hB9BA
`define CUBE_LUT_BB32 16'hB9BA
`define CUBE_LUT_BB33 16'hB9BB
`define CUBE_LUT_BB34 16'hB9BB
`define CUBE_LUT_BB35 16'hB9BC
`define CUBE_LUT_BB36 16'hB9BC
`define CUBE_LUT_BB37 16'hB9BD
`define CUBE_LUT_BB38 16'hB9BD
`define CUBE_LUT_BB39 16'hB9BE
`define CUBE_LUT_BB3A 16'hB9BE
`define CUBE_LUT_BB3B 16'hB9BF
`define CUBE_LUT_BB3C 16'hB9BF
`define CUBE_LUT_BB3D 16'hB9C0
`define CUBE_LUT_BB3E 16'hB9C0
`define CUBE_LUT_BB3F 16'hB9C1
`define CUBE_LUT_BB40 16'hB9C1
`define CUBE_LUT_BB41 16'hB9C2
`define CUBE_LUT_BB42 16'hB9C2
`define CUBE_LUT_BB43 16'hB9C3
`define CUBE_LUT_BB44 16'hB9C3
`define CUBE_LUT_BB45 16'hB9C4
`define CUBE_LUT_BB46 16'hB9C4
`define CUBE_LUT_BB47 16'hB9C5
`define CUBE_LUT_BB48 16'hB9C5
`define CUBE_LUT_BB49 16'hB9C6
`define CUBE_LUT_BB4A 16'hB9C6
`define CUBE_LUT_BB4B 16'hB9C6
`define CUBE_LUT_BB4C 16'hB9C7
`define CUBE_LUT_BB4D 16'hB9C7
`define CUBE_LUT_BB4E 16'hB9C8
`define CUBE_LUT_BB4F 16'hB9C8
`define CUBE_LUT_BB50 16'hB9C9
`define CUBE_LUT_BB51 16'hB9C9
`define CUBE_LUT_BB52 16'hB9CA
`define CUBE_LUT_BB53 16'hB9CA
`define CUBE_LUT_BB54 16'hB9CB
`define CUBE_LUT_BB55 16'hB9CB
`define CUBE_LUT_BB56 16'hB9CC
`define CUBE_LUT_BB57 16'hB9CC
`define CUBE_LUT_BB58 16'hB9CD
`define CUBE_LUT_BB59 16'hB9CD
`define CUBE_LUT_BB5A 16'hB9CE
`define CUBE_LUT_BB5B 16'hB9CE
`define CUBE_LUT_BB5C 16'hB9CF
`define CUBE_LUT_BB5D 16'hB9CF
`define CUBE_LUT_BB5E 16'hB9D0
`define CUBE_LUT_BB5F 16'hB9D0
`define CUBE_LUT_BB60 16'hB9D0
`define CUBE_LUT_BB61 16'hB9D1
`define CUBE_LUT_BB62 16'hB9D1
`define CUBE_LUT_BB63 16'hB9D2
`define CUBE_LUT_BB64 16'hB9D2
`define CUBE_LUT_BB65 16'hB9D3
`define CUBE_LUT_BB66 16'hB9D3
`define CUBE_LUT_BB67 16'hB9D4
`define CUBE_LUT_BB68 16'hB9D4
`define CUBE_LUT_BB69 16'hB9D5
`define CUBE_LUT_BB6A 16'hB9D5
`define CUBE_LUT_BB6B 16'hB9D6
`define CUBE_LUT_BB6C 16'hB9D6
`define CUBE_LUT_BB6D 16'hB9D7
`define CUBE_LUT_BB6E 16'hB9D7
`define CUBE_LUT_BB6F 16'hB9D7
`define CUBE_LUT_BB70 16'hB9D8
`define CUBE_LUT_BB71 16'hB9D8
`define CUBE_LUT_BB72 16'hB9D9
`define CUBE_LUT_BB73 16'hB9D9
`define CUBE_LUT_BB74 16'hB9DA
`define CUBE_LUT_BB75 16'hB9DA
`define CUBE_LUT_BB76 16'hB9DB
`define CUBE_LUT_BB77 16'hB9DB
`define CUBE_LUT_BB78 16'hB9DC
`define CUBE_LUT_BB79 16'hB9DC
`define CUBE_LUT_BB7A 16'hB9DD
`define CUBE_LUT_BB7B 16'hB9DD
`define CUBE_LUT_BB7C 16'hB9DE
`define CUBE_LUT_BB7D 16'hB9DE
`define CUBE_LUT_BB7E 16'hB9DE
`define CUBE_LUT_BB7F 16'hB9DF
`define CUBE_LUT_BB80 16'hB9DF
`define CUBE_LUT_BB81 16'hB9E0
`define CUBE_LUT_BB82 16'hB9E0
`define CUBE_LUT_BB83 16'hB9E1
`define CUBE_LUT_BB84 16'hB9E1
`define CUBE_LUT_BB85 16'hB9E2
`define CUBE_LUT_BB86 16'hB9E2
`define CUBE_LUT_BB87 16'hB9E3
`define CUBE_LUT_BB88 16'hB9E3
`define CUBE_LUT_BB89 16'hB9E4
`define CUBE_LUT_BB8A 16'hB9E4
`define CUBE_LUT_BB8B 16'hB9E4
`define CUBE_LUT_BB8C 16'hB9E5
`define CUBE_LUT_BB8D 16'hB9E5
`define CUBE_LUT_BB8E 16'hB9E6
`define CUBE_LUT_BB8F 16'hB9E6
`define CUBE_LUT_BB90 16'hB9E7
`define CUBE_LUT_BB91 16'hB9E7
`define CUBE_LUT_BB92 16'hB9E8
`define CUBE_LUT_BB93 16'hB9E8
`define CUBE_LUT_BB94 16'hB9E9
`define CUBE_LUT_BB95 16'hB9E9
`define CUBE_LUT_BB96 16'hB9E9
`define CUBE_LUT_BB97 16'hB9EA
`define CUBE_LUT_BB98 16'hB9EA
`define CUBE_LUT_BB99 16'hB9EB
`define CUBE_LUT_BB9A 16'hB9EB
`define CUBE_LUT_BB9B 16'hB9EC
`define CUBE_LUT_BB9C 16'hB9EC
`define CUBE_LUT_BB9D 16'hB9ED
`define CUBE_LUT_BB9E 16'hB9ED
`define CUBE_LUT_BB9F 16'hB9EE
`define CUBE_LUT_BBA0 16'hB9EE
`define CUBE_LUT_BBA1 16'hB9EE
`define CUBE_LUT_BBA2 16'hB9EF
`define CUBE_LUT_BBA3 16'hB9EF
`define CUBE_LUT_BBA4 16'hB9F0
`define CUBE_LUT_BBA5 16'hB9F0
`define CUBE_LUT_BBA6 16'hB9F1
`define CUBE_LUT_BBA7 16'hB9F1
`define CUBE_LUT_BBA8 16'hB9F2
`define CUBE_LUT_BBA9 16'hB9F2
`define CUBE_LUT_BBAA 16'hB9F2
`define CUBE_LUT_BBAB 16'hB9F3
`define CUBE_LUT_BBAC 16'hB9F3
`define CUBE_LUT_BBAD 16'hB9F4
`define CUBE_LUT_BBAE 16'hB9F4
`define CUBE_LUT_BBAF 16'hB9F5
`define CUBE_LUT_BBB0 16'hB9F5
`define CUBE_LUT_BBB1 16'hB9F6
`define CUBE_LUT_BBB2 16'hB9F6
`define CUBE_LUT_BBB3 16'hB9F6
`define CUBE_LUT_BBB4 16'hB9F7
`define CUBE_LUT_BBB5 16'hB9F7
`define CUBE_LUT_BBB6 16'hB9F8
`define CUBE_LUT_BBB7 16'hB9F8
`define CUBE_LUT_BBB8 16'hB9F9
`define CUBE_LUT_BBB9 16'hB9F9
`define CUBE_LUT_BBBA 16'hB9FA
`define CUBE_LUT_BBBB 16'hB9FA
`define CUBE_LUT_BBBC 16'hB9FA
`define CUBE_LUT_BBBD 16'hB9FB
`define CUBE_LUT_BBBE 16'hB9FB
`define CUBE_LUT_BBBF 16'hB9FC
`define CUBE_LUT_BBC0 16'hB9FC
`define CUBE_LUT_BBC1 16'hB9FD
`define CUBE_LUT_BBC2 16'hB9FD
`define CUBE_LUT_BBC3 16'hB9FE
`define CUBE_LUT_BBC4 16'hB9FE
`define CUBE_LUT_BBC5 16'hB9FE
`define CUBE_LUT_BBC6 16'hB9FF
`define CUBE_LUT_BBC7 16'hB9FF
`define CUBE_LUT_BBC8 16'hBA00
`define CUBE_LUT_BBC9 16'hBA00
`define CUBE_LUT_BBCA 16'hBA01
`define CUBE_LUT_BBCB 16'hBA01
`define CUBE_LUT_BBCC 16'hBA01
`define CUBE_LUT_BBCD 16'hBA02
`define CUBE_LUT_BBCE 16'hBA02
`define CUBE_LUT_BBCF 16'hBA03
`define CUBE_LUT_BBD0 16'hBA03
`define CUBE_LUT_BBD1 16'hBA04
`define CUBE_LUT_BBD2 16'hBA04
`define CUBE_LUT_BBD3 16'hBA05
`define CUBE_LUT_BBD4 16'hBA05
`define CUBE_LUT_BBD5 16'hBA05
`define CUBE_LUT_BBD6 16'hBA06
`define CUBE_LUT_BBD7 16'hBA06
`define CUBE_LUT_BBD8 16'hBA07
`define CUBE_LUT_BBD9 16'hBA07
`define CUBE_LUT_BBDA 16'hBA08
`define CUBE_LUT_BBDB 16'hBA08
`define CUBE_LUT_BBDC 16'hBA08
`define CUBE_LUT_BBDD 16'hBA09
`define CUBE_LUT_BBDE 16'hBA09
`define CUBE_LUT_BBDF 16'hBA0A
`define CUBE_LUT_BBE0 16'hBA0A
`define CUBE_LUT_BBE1 16'hBA0B
`define CUBE_LUT_BBE2 16'hBA0B
`define CUBE_LUT_BBE3 16'hBA0B
`define CUBE_LUT_BBE4 16'hBA0C
`define CUBE_LUT_BBE5 16'hBA0C
`define CUBE_LUT_BBE6 16'hBA0D
`define CUBE_LUT_BBE7 16'hBA0D
`define CUBE_LUT_BBE8 16'hBA0E
`define CUBE_LUT_BBE9 16'hBA0E
`define CUBE_LUT_BBEA 16'hBA0E
`define CUBE_LUT_BBEB 16'hBA0F
`define CUBE_LUT_BBEC 16'hBA0F
`define CUBE_LUT_BBED 16'hBA10
`define CUBE_LUT_BBEE 16'hBA10
`define CUBE_LUT_BBEF 16'hBA11
`define CUBE_LUT_BBF0 16'hBA11
`define CUBE_LUT_BBF1 16'hBA11
`define CUBE_LUT_BBF2 16'hBA12
`define CUBE_LUT_BBF3 16'hBA12
`define CUBE_LUT_BBF4 16'hBA13
`define CUBE_LUT_BBF5 16'hBA13
`define CUBE_LUT_BBF6 16'hBA14
`define CUBE_LUT_BBF7 16'hBA14
`define CUBE_LUT_BBF8 16'hBA14
`define CUBE_LUT_BBF9 16'hBA15
`define CUBE_LUT_BBFA 16'hBA15
`define CUBE_LUT_BBFB 16'hBA16
`define CUBE_LUT_BBFC 16'hBA16
`define CUBE_LUT_BBFD 16'hBA16
`define CUBE_LUT_BBFE 16'hBA17
`define CUBE_LUT_BBFF 16'hBA17
`define CUBE_LUT_BC00 16'hBA18
`define CUBE_LUT_BC01 16'hBA19
`define CUBE_LUT_BC02 16'hBA19
`define CUBE_LUT_BC03 16'hBA1A
`define CUBE_LUT_BC04 16'hBA1B
`define CUBE_LUT_BC05 16'hBA1C
`define CUBE_LUT_BC06 16'hBA1D
`define CUBE_LUT_BC07 16'hBA1E
`define CUBE_LUT_BC08 16'hBA1E
`define CUBE_LUT_BC09 16'hBA1F
`define CUBE_LUT_BC0A 16'hBA20
`define CUBE_LUT_BC0B 16'hBA21
`define CUBE_LUT_BC0C 16'hBA22
`define CUBE_LUT_BC0D 16'hBA23
`define CUBE_LUT_BC0E 16'hBA23
`define CUBE_LUT_BC0F 16'hBA24
`define CUBE_LUT_BC10 16'hBA25
`define CUBE_LUT_BC11 16'hBA26
`define CUBE_LUT_BC12 16'hBA27
`define CUBE_LUT_BC13 16'hBA27
`define CUBE_LUT_BC14 16'hBA28
`define CUBE_LUT_BC15 16'hBA29
`define CUBE_LUT_BC16 16'hBA2A
`define CUBE_LUT_BC17 16'hBA2B
`define CUBE_LUT_BC18 16'hBA2C
`define CUBE_LUT_BC19 16'hBA2C
`define CUBE_LUT_BC1A 16'hBA2D
`define CUBE_LUT_BC1B 16'hBA2E
`define CUBE_LUT_BC1C 16'hBA2F
`define CUBE_LUT_BC1D 16'hBA30
`define CUBE_LUT_BC1E 16'hBA30
`define CUBE_LUT_BC1F 16'hBA31
`define CUBE_LUT_BC20 16'hBA32
`define CUBE_LUT_BC21 16'hBA33
`define CUBE_LUT_BC22 16'hBA34
`define CUBE_LUT_BC23 16'hBA34
`define CUBE_LUT_BC24 16'hBA35
`define CUBE_LUT_BC25 16'hBA36
`define CUBE_LUT_BC26 16'hBA37
`define CUBE_LUT_BC27 16'hBA38
`define CUBE_LUT_BC28 16'hBA38
`define CUBE_LUT_BC29 16'hBA39
`define CUBE_LUT_BC2A 16'hBA3A
`define CUBE_LUT_BC2B 16'hBA3B
`define CUBE_LUT_BC2C 16'hBA3C
`define CUBE_LUT_BC2D 16'hBA3C
`define CUBE_LUT_BC2E 16'hBA3D
`define CUBE_LUT_BC2F 16'hBA3E
`define CUBE_LUT_BC30 16'hBA3F
`define CUBE_LUT_BC31 16'hBA3F
`define CUBE_LUT_BC32 16'hBA40
`define CUBE_LUT_BC33 16'hBA41
`define CUBE_LUT_BC34 16'hBA42
`define CUBE_LUT_BC35 16'hBA43
`define CUBE_LUT_BC36 16'hBA43
`define CUBE_LUT_BC37 16'hBA44
`define CUBE_LUT_BC38 16'hBA45
`define CUBE_LUT_BC39 16'hBA46
`define CUBE_LUT_BC3A 16'hBA46
`define CUBE_LUT_BC3B 16'hBA47
`define CUBE_LUT_BC3C 16'hBA48
`define CUBE_LUT_BC3D 16'hBA49
`define CUBE_LUT_BC3E 16'hBA49
`define CUBE_LUT_BC3F 16'hBA4A
`define CUBE_LUT_BC40 16'hBA4B
`define CUBE_LUT_BC41 16'hBA4C
`define CUBE_LUT_BC42 16'hBA4D
`define CUBE_LUT_BC43 16'hBA4D
`define CUBE_LUT_BC44 16'hBA4E
`define CUBE_LUT_BC45 16'hBA4F
`define CUBE_LUT_BC46 16'hBA50
`define CUBE_LUT_BC47 16'hBA50
`define CUBE_LUT_BC48 16'hBA51
`define CUBE_LUT_BC49 16'hBA52
`define CUBE_LUT_BC4A 16'hBA53
`define CUBE_LUT_BC4B 16'hBA53
`define CUBE_LUT_BC4C 16'hBA54
`define CUBE_LUT_BC4D 16'hBA55
`define CUBE_LUT_BC4E 16'hBA56
`define CUBE_LUT_BC4F 16'hBA56
`define CUBE_LUT_BC50 16'hBA57
`define CUBE_LUT_BC51 16'hBA58
`define CUBE_LUT_BC52 16'hBA59
`define CUBE_LUT_BC53 16'hBA59
`define CUBE_LUT_BC54 16'hBA5A
`define CUBE_LUT_BC55 16'hBA5B
`define CUBE_LUT_BC56 16'hBA5B
`define CUBE_LUT_BC57 16'hBA5C
`define CUBE_LUT_BC58 16'hBA5D
`define CUBE_LUT_BC59 16'hBA5E
`define CUBE_LUT_BC5A 16'hBA5E
`define CUBE_LUT_BC5B 16'hBA5F
`define CUBE_LUT_BC5C 16'hBA60
`define CUBE_LUT_BC5D 16'hBA61
`define CUBE_LUT_BC5E 16'hBA61
`define CUBE_LUT_BC5F 16'hBA62
`define CUBE_LUT_BC60 16'hBA63
`define CUBE_LUT_BC61 16'hBA64
`define CUBE_LUT_BC62 16'hBA64
`define CUBE_LUT_BC63 16'hBA65
`define CUBE_LUT_BC64 16'hBA66
`define CUBE_LUT_BC65 16'hBA66
`define CUBE_LUT_BC66 16'hBA67
`define CUBE_LUT_BC67 16'hBA68
`define CUBE_LUT_BC68 16'hBA69
`define CUBE_LUT_BC69 16'hBA69
`define CUBE_LUT_BC6A 16'hBA6A
`define CUBE_LUT_BC6B 16'hBA6B
`define CUBE_LUT_BC6C 16'hBA6B
`define CUBE_LUT_BC6D 16'hBA6C
`define CUBE_LUT_BC6E 16'hBA6D
`define CUBE_LUT_BC6F 16'hBA6E
`define CUBE_LUT_BC70 16'hBA6E
`define CUBE_LUT_BC71 16'hBA6F
`define CUBE_LUT_BC72 16'hBA70
`define CUBE_LUT_BC73 16'hBA70
`define CUBE_LUT_BC74 16'hBA71
`define CUBE_LUT_BC75 16'hBA72
`define CUBE_LUT_BC76 16'hBA72
`define CUBE_LUT_BC77 16'hBA73
`define CUBE_LUT_BC78 16'hBA74
`define CUBE_LUT_BC79 16'hBA75
`define CUBE_LUT_BC7A 16'hBA75
`define CUBE_LUT_BC7B 16'hBA76
`define CUBE_LUT_BC7C 16'hBA77
`define CUBE_LUT_BC7D 16'hBA77
`define CUBE_LUT_BC7E 16'hBA78
`define CUBE_LUT_BC7F 16'hBA79
`define CUBE_LUT_BC80 16'hBA79
`define CUBE_LUT_BC81 16'hBA7A
`define CUBE_LUT_BC82 16'hBA7B
`define CUBE_LUT_BC83 16'hBA7C
`define CUBE_LUT_BC84 16'hBA7C
`define CUBE_LUT_BC85 16'hBA7D
`define CUBE_LUT_BC86 16'hBA7E
`define CUBE_LUT_BC87 16'hBA7E
`define CUBE_LUT_BC88 16'hBA7F
`define CUBE_LUT_BC89 16'hBA80
`define CUBE_LUT_BC8A 16'hBA80
`define CUBE_LUT_BC8B 16'hBA81
`define CUBE_LUT_BC8C 16'hBA82
`define CUBE_LUT_BC8D 16'hBA82
`define CUBE_LUT_BC8E 16'hBA83
`define CUBE_LUT_BC8F 16'hBA84
`define CUBE_LUT_BC90 16'hBA84
`define CUBE_LUT_BC91 16'hBA85
`define CUBE_LUT_BC92 16'hBA86
`define CUBE_LUT_BC93 16'hBA86
`define CUBE_LUT_BC94 16'hBA87
`define CUBE_LUT_BC95 16'hBA88
`define CUBE_LUT_BC96 16'hBA88
`define CUBE_LUT_BC97 16'hBA89
`define CUBE_LUT_BC98 16'hBA8A
`define CUBE_LUT_BC99 16'hBA8A
`define CUBE_LUT_BC9A 16'hBA8B
`define CUBE_LUT_BC9B 16'hBA8C
`define CUBE_LUT_BC9C 16'hBA8C
`define CUBE_LUT_BC9D 16'hBA8D
`define CUBE_LUT_BC9E 16'hBA8E
`define CUBE_LUT_BC9F 16'hBA8E
`define CUBE_LUT_BCA0 16'hBA8F
`define CUBE_LUT_BCA1 16'hBA90
`define CUBE_LUT_BCA2 16'hBA90
`define CUBE_LUT_BCA3 16'hBA91
`define CUBE_LUT_BCA4 16'hBA92
`define CUBE_LUT_BCA5 16'hBA92
`define CUBE_LUT_BCA6 16'hBA93
`define CUBE_LUT_BCA7 16'hBA94
`define CUBE_LUT_BCA8 16'hBA94
`define CUBE_LUT_BCA9 16'hBA95
`define CUBE_LUT_BCAA 16'hBA95
`define CUBE_LUT_BCAB 16'hBA96
`define CUBE_LUT_BCAC 16'hBA97
`define CUBE_LUT_BCAD 16'hBA97
`define CUBE_LUT_BCAE 16'hBA98
`define CUBE_LUT_BCAF 16'hBA99
`define CUBE_LUT_BCB0 16'hBA99
`define CUBE_LUT_BCB1 16'hBA9A
`define CUBE_LUT_BCB2 16'hBA9B
`define CUBE_LUT_BCB3 16'hBA9B
`define CUBE_LUT_BCB4 16'hBA9C
`define CUBE_LUT_BCB5 16'hBA9D
`define CUBE_LUT_BCB6 16'hBA9D
`define CUBE_LUT_BCB7 16'hBA9E
`define CUBE_LUT_BCB8 16'hBA9E
`define CUBE_LUT_BCB9 16'hBA9F
`define CUBE_LUT_BCBA 16'hBAA0
`define CUBE_LUT_BCBB 16'hBAA0
`define CUBE_LUT_BCBC 16'hBAA1
`define CUBE_LUT_BCBD 16'hBAA2
`define CUBE_LUT_BCBE 16'hBAA2
`define CUBE_LUT_BCBF 16'hBAA3
`define CUBE_LUT_BCC0 16'hBAA3
`define CUBE_LUT_BCC1 16'hBAA4
`define CUBE_LUT_BCC2 16'hBAA5
`define CUBE_LUT_BCC3 16'hBAA5
`define CUBE_LUT_BCC4 16'hBAA6
`define CUBE_LUT_BCC5 16'hBAA7
`define CUBE_LUT_BCC6 16'hBAA7
`define CUBE_LUT_BCC7 16'hBAA8
`define CUBE_LUT_BCC8 16'hBAA8
`define CUBE_LUT_BCC9 16'hBAA9
`define CUBE_LUT_BCCA 16'hBAAA
`define CUBE_LUT_BCCB 16'hBAAA
`define CUBE_LUT_BCCC 16'hBAAB
`define CUBE_LUT_BCCD 16'hBAAB
`define CUBE_LUT_BCCE 16'hBAAC
`define CUBE_LUT_BCCF 16'hBAAD
`define CUBE_LUT_BCD0 16'hBAAD
`define CUBE_LUT_BCD1 16'hBAAE
`define CUBE_LUT_BCD2 16'hBAAE
`define CUBE_LUT_BCD3 16'hBAAF
`define CUBE_LUT_BCD4 16'hBAB0
`define CUBE_LUT_BCD5 16'hBAB0
`define CUBE_LUT_BCD6 16'hBAB1
`define CUBE_LUT_BCD7 16'hBAB1
`define CUBE_LUT_BCD8 16'hBAB2
`define CUBE_LUT_BCD9 16'hBAB3
`define CUBE_LUT_BCDA 16'hBAB3
`define CUBE_LUT_BCDB 16'hBAB4
`define CUBE_LUT_BCDC 16'hBAB4
`define CUBE_LUT_BCDD 16'hBAB5
`define CUBE_LUT_BCDE 16'hBAB6
`define CUBE_LUT_BCDF 16'hBAB6
`define CUBE_LUT_BCE0 16'hBAB7
`define CUBE_LUT_BCE1 16'hBAB7
`define CUBE_LUT_BCE2 16'hBAB8
`define CUBE_LUT_BCE3 16'hBAB9
`define CUBE_LUT_BCE4 16'hBAB9
`define CUBE_LUT_BCE5 16'hBABA
`define CUBE_LUT_BCE6 16'hBABA
`define CUBE_LUT_BCE7 16'hBABB
`define CUBE_LUT_BCE8 16'hBABC
`define CUBE_LUT_BCE9 16'hBABC
`define CUBE_LUT_BCEA 16'hBABD
`define CUBE_LUT_BCEB 16'hBABD
`define CUBE_LUT_BCEC 16'hBABE
`define CUBE_LUT_BCED 16'hBABE
`define CUBE_LUT_BCEE 16'hBABF
`define CUBE_LUT_BCEF 16'hBAC0
`define CUBE_LUT_BCF0 16'hBAC0
`define CUBE_LUT_BCF1 16'hBAC1
`define CUBE_LUT_BCF2 16'hBAC1
`define CUBE_LUT_BCF3 16'hBAC2
`define CUBE_LUT_BCF4 16'hBAC2
`define CUBE_LUT_BCF5 16'hBAC3
`define CUBE_LUT_BCF6 16'hBAC4
`define CUBE_LUT_BCF7 16'hBAC4
`define CUBE_LUT_BCF8 16'hBAC5
`define CUBE_LUT_BCF9 16'hBAC5
`define CUBE_LUT_BCFA 16'hBAC6
`define CUBE_LUT_BCFB 16'hBAC6
`define CUBE_LUT_BCFC 16'hBAC7
`define CUBE_LUT_BCFD 16'hBAC8
`define CUBE_LUT_BCFE 16'hBAC8
`define CUBE_LUT_BCFF 16'hBAC9
`define CUBE_LUT_BD00 16'hBAC9
`define CUBE_LUT_BD01 16'hBACA
`define CUBE_LUT_BD02 16'hBACA
`define CUBE_LUT_BD03 16'hBACB
`define CUBE_LUT_BD04 16'hBACC
`define CUBE_LUT_BD05 16'hBACC
`define CUBE_LUT_BD06 16'hBACD
`define CUBE_LUT_BD07 16'hBACD
`define CUBE_LUT_BD08 16'hBACE
`define CUBE_LUT_BD09 16'hBACE
`define CUBE_LUT_BD0A 16'hBACF
`define CUBE_LUT_BD0B 16'hBACF
`define CUBE_LUT_BD0C 16'hBAD0
`define CUBE_LUT_BD0D 16'hBAD0
`define CUBE_LUT_BD0E 16'hBAD1
`define CUBE_LUT_BD0F 16'hBAD2
`define CUBE_LUT_BD10 16'hBAD2
`define CUBE_LUT_BD11 16'hBAD3
`define CUBE_LUT_BD12 16'hBAD3
`define CUBE_LUT_BD13 16'hBAD4
`define CUBE_LUT_BD14 16'hBAD4
`define CUBE_LUT_BD15 16'hBAD5
`define CUBE_LUT_BD16 16'hBAD5
`define CUBE_LUT_BD17 16'hBAD6
`define CUBE_LUT_BD18 16'hBAD6
`define CUBE_LUT_BD19 16'hBAD7
`define CUBE_LUT_BD1A 16'hBAD8
`define CUBE_LUT_BD1B 16'hBAD8
`define CUBE_LUT_BD1C 16'hBAD9
`define CUBE_LUT_BD1D 16'hBAD9
`define CUBE_LUT_BD1E 16'hBADA
`define CUBE_LUT_BD1F 16'hBADA
`define CUBE_LUT_BD20 16'hBADB
`define CUBE_LUT_BD21 16'hBADB
`define CUBE_LUT_BD22 16'hBADC
`define CUBE_LUT_BD23 16'hBADC
`define CUBE_LUT_BD24 16'hBADD
`define CUBE_LUT_BD25 16'hBADD
`define CUBE_LUT_BD26 16'hBADE
`define CUBE_LUT_BD27 16'hBADE
`define CUBE_LUT_BD28 16'hBADF
`define CUBE_LUT_BD29 16'hBAE0
`define CUBE_LUT_BD2A 16'hBAE0
`define CUBE_LUT_BD2B 16'hBAE1
`define CUBE_LUT_BD2C 16'hBAE1
`define CUBE_LUT_BD2D 16'hBAE2
`define CUBE_LUT_BD2E 16'hBAE2
`define CUBE_LUT_BD2F 16'hBAE3
`define CUBE_LUT_BD30 16'hBAE3
`define CUBE_LUT_BD31 16'hBAE4
`define CUBE_LUT_BD32 16'hBAE4
`define CUBE_LUT_BD33 16'hBAE5
`define CUBE_LUT_BD34 16'hBAE5
`define CUBE_LUT_BD35 16'hBAE6
`define CUBE_LUT_BD36 16'hBAE6
`define CUBE_LUT_BD37 16'hBAE7
`define CUBE_LUT_BD38 16'hBAE7
`define CUBE_LUT_BD39 16'hBAE8
`define CUBE_LUT_BD3A 16'hBAE8
`define CUBE_LUT_BD3B 16'hBAE9
`define CUBE_LUT_BD3C 16'hBAE9
`define CUBE_LUT_BD3D 16'hBAEA
`define CUBE_LUT_BD3E 16'hBAEA
`define CUBE_LUT_BD3F 16'hBAEB
`define CUBE_LUT_BD40 16'hBAEB
`define CUBE_LUT_BD41 16'hBAEC
`define CUBE_LUT_BD42 16'hBAEC
`define CUBE_LUT_BD43 16'hBAED
`define CUBE_LUT_BD44 16'hBAED
`define CUBE_LUT_BD45 16'hBAEE
`define CUBE_LUT_BD46 16'hBAEE
`define CUBE_LUT_BD47 16'hBAEF
`define CUBE_LUT_BD48 16'hBAEF
`define CUBE_LUT_BD49 16'hBAF0
`define CUBE_LUT_BD4A 16'hBAF0
`define CUBE_LUT_BD4B 16'hBAF1
`define CUBE_LUT_BD4C 16'hBAF1
`define CUBE_LUT_BD4D 16'hBAF2
`define CUBE_LUT_BD4E 16'hBAF2
`define CUBE_LUT_BD4F 16'hBAF3
`define CUBE_LUT_BD50 16'hBAF3
`define CUBE_LUT_BD51 16'hBAF4
`define CUBE_LUT_BD52 16'hBAF4
`define CUBE_LUT_BD53 16'hBAF5
`define CUBE_LUT_BD54 16'hBAF5
`define CUBE_LUT_BD55 16'hBAF6
`define CUBE_LUT_BD56 16'hBAF6
`define CUBE_LUT_BD57 16'hBAF7
`define CUBE_LUT_BD58 16'hBAF7
`define CUBE_LUT_BD59 16'hBAF8
`define CUBE_LUT_BD5A 16'hBAF8
`define CUBE_LUT_BD5B 16'hBAF9
`define CUBE_LUT_BD5C 16'hBAF9
`define CUBE_LUT_BD5D 16'hBAFA
`define CUBE_LUT_BD5E 16'hBAFA
`define CUBE_LUT_BD5F 16'hBAFB
`define CUBE_LUT_BD60 16'hBAFB
`define CUBE_LUT_BD61 16'hBAFC
`define CUBE_LUT_BD62 16'hBAFC
`define CUBE_LUT_BD63 16'hBAFC
`define CUBE_LUT_BD64 16'hBAFD
`define CUBE_LUT_BD65 16'hBAFD
`define CUBE_LUT_BD66 16'hBAFE
`define CUBE_LUT_BD67 16'hBAFE
`define CUBE_LUT_BD68 16'hBAFF
`define CUBE_LUT_BD69 16'hBAFF
`define CUBE_LUT_BD6A 16'hBB00
`define CUBE_LUT_BD6B 16'hBB00
`define CUBE_LUT_BD6C 16'hBB01
`define CUBE_LUT_BD6D 16'hBB01
`define CUBE_LUT_BD6E 16'hBB02
`define CUBE_LUT_BD6F 16'hBB02
`define CUBE_LUT_BD70 16'hBB03
`define CUBE_LUT_BD71 16'hBB03
`define CUBE_LUT_BD72 16'hBB03
`define CUBE_LUT_BD73 16'hBB04
`define CUBE_LUT_BD74 16'hBB04
`define CUBE_LUT_BD75 16'hBB05
`define CUBE_LUT_BD76 16'hBB05
`define CUBE_LUT_BD77 16'hBB06
`define CUBE_LUT_BD78 16'hBB06
`define CUBE_LUT_BD79 16'hBB07
`define CUBE_LUT_BD7A 16'hBB07
`define CUBE_LUT_BD7B 16'hBB08
`define CUBE_LUT_BD7C 16'hBB08
`define CUBE_LUT_BD7D 16'hBB09
`define CUBE_LUT_BD7E 16'hBB09
`define CUBE_LUT_BD7F 16'hBB09
`define CUBE_LUT_BD80 16'hBB0A
`define CUBE_LUT_BD81 16'hBB0A
`define CUBE_LUT_BD82 16'hBB0B
`define CUBE_LUT_BD83 16'hBB0B
`define CUBE_LUT_BD84 16'hBB0C
`define CUBE_LUT_BD85 16'hBB0C
`define CUBE_LUT_BD86 16'hBB0D
`define CUBE_LUT_BD87 16'hBB0D
`define CUBE_LUT_BD88 16'hBB0D
`define CUBE_LUT_BD89 16'hBB0E
`define CUBE_LUT_BD8A 16'hBB0E
`define CUBE_LUT_BD8B 16'hBB0F
`define CUBE_LUT_BD8C 16'hBB0F
`define CUBE_LUT_BD8D 16'hBB10
`define CUBE_LUT_BD8E 16'hBB10
`define CUBE_LUT_BD8F 16'hBB11
`define CUBE_LUT_BD90 16'hBB11
`define CUBE_LUT_BD91 16'hBB11
`define CUBE_LUT_BD92 16'hBB12
`define CUBE_LUT_BD93 16'hBB12
`define CUBE_LUT_BD94 16'hBB13
`define CUBE_LUT_BD95 16'hBB13
`define CUBE_LUT_BD96 16'hBB14
`define CUBE_LUT_BD97 16'hBB14
`define CUBE_LUT_BD98 16'hBB15
`define CUBE_LUT_BD99 16'hBB15
`define CUBE_LUT_BD9A 16'hBB15
`define CUBE_LUT_BD9B 16'hBB16
`define CUBE_LUT_BD9C 16'hBB16
`define CUBE_LUT_BD9D 16'hBB17
`define CUBE_LUT_BD9E 16'hBB17
`define CUBE_LUT_BD9F 16'hBB18
`define CUBE_LUT_BDA0 16'hBB18
`define CUBE_LUT_BDA1 16'hBB18
`define CUBE_LUT_BDA2 16'hBB19
`define CUBE_LUT_BDA3 16'hBB19
`define CUBE_LUT_BDA4 16'hBB1A
`define CUBE_LUT_BDA5 16'hBB1A
`define CUBE_LUT_BDA6 16'hBB1B
`define CUBE_LUT_BDA7 16'hBB1B
`define CUBE_LUT_BDA8 16'hBB1B
`define CUBE_LUT_BDA9 16'hBB1C
`define CUBE_LUT_BDAA 16'hBB1C
`define CUBE_LUT_BDAB 16'hBB1D
`define CUBE_LUT_BDAC 16'hBB1D
`define CUBE_LUT_BDAD 16'hBB1D
`define CUBE_LUT_BDAE 16'hBB1E
`define CUBE_LUT_BDAF 16'hBB1E
`define CUBE_LUT_BDB0 16'hBB1F
`define CUBE_LUT_BDB1 16'hBB1F
`define CUBE_LUT_BDB2 16'hBB20
`define CUBE_LUT_BDB3 16'hBB20
`define CUBE_LUT_BDB4 16'hBB20
`define CUBE_LUT_BDB5 16'hBB21
`define CUBE_LUT_BDB6 16'hBB21
`define CUBE_LUT_BDB7 16'hBB22
`define CUBE_LUT_BDB8 16'hBB22
`define CUBE_LUT_BDB9 16'hBB22
`define CUBE_LUT_BDBA 16'hBB23
`define CUBE_LUT_BDBB 16'hBB23
`define CUBE_LUT_BDBC 16'hBB24
`define CUBE_LUT_BDBD 16'hBB24
`define CUBE_LUT_BDBE 16'hBB24
`define CUBE_LUT_BDBF 16'hBB25
`define CUBE_LUT_BDC0 16'hBB25
`define CUBE_LUT_BDC1 16'hBB26
`define CUBE_LUT_BDC2 16'hBB26
`define CUBE_LUT_BDC3 16'hBB26
`define CUBE_LUT_BDC4 16'hBB27
`define CUBE_LUT_BDC5 16'hBB27
`define CUBE_LUT_BDC6 16'hBB28
`define CUBE_LUT_BDC7 16'hBB28
`define CUBE_LUT_BDC8 16'hBB28
`define CUBE_LUT_BDC9 16'hBB29
`define CUBE_LUT_BDCA 16'hBB29
`define CUBE_LUT_BDCB 16'hBB2A
`define CUBE_LUT_BDCC 16'hBB2A
`define CUBE_LUT_BDCD 16'hBB2A
`define CUBE_LUT_BDCE 16'hBB2B
`define CUBE_LUT_BDCF 16'hBB2B
`define CUBE_LUT_BDD0 16'hBB2C
`define CUBE_LUT_BDD1 16'hBB2C
`define CUBE_LUT_BDD2 16'hBB2C
`define CUBE_LUT_BDD3 16'hBB2D
`define CUBE_LUT_BDD4 16'hBB2D
`define CUBE_LUT_BDD5 16'hBB2E
`define CUBE_LUT_BDD6 16'hBB2E
`define CUBE_LUT_BDD7 16'hBB2E
`define CUBE_LUT_BDD8 16'hBB2F
`define CUBE_LUT_BDD9 16'hBB2F
`define CUBE_LUT_BDDA 16'hBB30
`define CUBE_LUT_BDDB 16'hBB30
`define CUBE_LUT_BDDC 16'hBB30
`define CUBE_LUT_BDDD 16'hBB31
`define CUBE_LUT_BDDE 16'hBB31
`define CUBE_LUT_BDDF 16'hBB31
`define CUBE_LUT_BDE0 16'hBB32
`define CUBE_LUT_BDE1 16'hBB32
`define CUBE_LUT_BDE2 16'hBB33
`define CUBE_LUT_BDE3 16'hBB33
`define CUBE_LUT_BDE4 16'hBB33
`define CUBE_LUT_BDE5 16'hBB34
`define CUBE_LUT_BDE6 16'hBB34
`define CUBE_LUT_BDE7 16'hBB35
`define CUBE_LUT_BDE8 16'hBB35
`define CUBE_LUT_BDE9 16'hBB35
`define CUBE_LUT_BDEA 16'hBB36
`define CUBE_LUT_BDEB 16'hBB36
`define CUBE_LUT_BDEC 16'hBB36
`define CUBE_LUT_BDED 16'hBB37
`define CUBE_LUT_BDEE 16'hBB37
`define CUBE_LUT_BDEF 16'hBB38
`define CUBE_LUT_BDF0 16'hBB38
`define CUBE_LUT_BDF1 16'hBB38
`define CUBE_LUT_BDF2 16'hBB39
`define CUBE_LUT_BDF3 16'hBB39
`define CUBE_LUT_BDF4 16'hBB39
`define CUBE_LUT_BDF5 16'hBB3A
`define CUBE_LUT_BDF6 16'hBB3A
`define CUBE_LUT_BDF7 16'hBB3A
`define CUBE_LUT_BDF8 16'hBB3B
`define CUBE_LUT_BDF9 16'hBB3B
`define CUBE_LUT_BDFA 16'hBB3C
`define CUBE_LUT_BDFB 16'hBB3C
`define CUBE_LUT_BDFC 16'hBB3C
`define CUBE_LUT_BDFD 16'hBB3D
`define CUBE_LUT_BDFE 16'hBB3D
`define CUBE_LUT_BDFF 16'hBB3D
`define CUBE_LUT_BE00 16'hBB3E
`define CUBE_LUT_BE01 16'hBB3E
`define CUBE_LUT_BE02 16'hBB3E
`define CUBE_LUT_BE03 16'hBB3F
`define CUBE_LUT_BE04 16'hBB3F
`define CUBE_LUT_BE05 16'hBB40
`define CUBE_LUT_BE06 16'hBB40
`define CUBE_LUT_BE07 16'hBB40
`define CUBE_LUT_BE08 16'hBB41
`define CUBE_LUT_BE09 16'hBB41
`define CUBE_LUT_BE0A 16'hBB41
`define CUBE_LUT_BE0B 16'hBB42
`define CUBE_LUT_BE0C 16'hBB42
`define CUBE_LUT_BE0D 16'hBB42
`define CUBE_LUT_BE0E 16'hBB43
`define CUBE_LUT_BE0F 16'hBB43
`define CUBE_LUT_BE10 16'hBB43
`define CUBE_LUT_BE11 16'hBB44
`define CUBE_LUT_BE12 16'hBB44
`define CUBE_LUT_BE13 16'hBB44
`define CUBE_LUT_BE14 16'hBB45
`define CUBE_LUT_BE15 16'hBB45
`define CUBE_LUT_BE16 16'hBB46
`define CUBE_LUT_BE17 16'hBB46
`define CUBE_LUT_BE18 16'hBB46
`define CUBE_LUT_BE19 16'hBB47
`define CUBE_LUT_BE1A 16'hBB47
`define CUBE_LUT_BE1B 16'hBB47
`define CUBE_LUT_BE1C 16'hBB48
`define CUBE_LUT_BE1D 16'hBB48
`define CUBE_LUT_BE1E 16'hBB48
`define CUBE_LUT_BE1F 16'hBB49
`define CUBE_LUT_BE20 16'hBB49
`define CUBE_LUT_BE21 16'hBB49
`define CUBE_LUT_BE22 16'hBB4A
`define CUBE_LUT_BE23 16'hBB4A
`define CUBE_LUT_BE24 16'hBB4A
`define CUBE_LUT_BE25 16'hBB4B
`define CUBE_LUT_BE26 16'hBB4B
`define CUBE_LUT_BE27 16'hBB4B
`define CUBE_LUT_BE28 16'hBB4C
`define CUBE_LUT_BE29 16'hBB4C
`define CUBE_LUT_BE2A 16'hBB4C
`define CUBE_LUT_BE2B 16'hBB4D
`define CUBE_LUT_BE2C 16'hBB4D
`define CUBE_LUT_BE2D 16'hBB4D
`define CUBE_LUT_BE2E 16'hBB4E
`define CUBE_LUT_BE2F 16'hBB4E
`define CUBE_LUT_BE30 16'hBB4E
`define CUBE_LUT_BE31 16'hBB4F
`define CUBE_LUT_BE32 16'hBB4F
`define CUBE_LUT_BE33 16'hBB4F
`define CUBE_LUT_BE34 16'hBB50
`define CUBE_LUT_BE35 16'hBB50
`define CUBE_LUT_BE36 16'hBB50
`define CUBE_LUT_BE37 16'hBB51
`define CUBE_LUT_BE38 16'hBB51
`define CUBE_LUT_BE39 16'hBB51
`define CUBE_LUT_BE3A 16'hBB52
`define CUBE_LUT_BE3B 16'hBB52
`define CUBE_LUT_BE3C 16'hBB52
`define CUBE_LUT_BE3D 16'hBB53
`define CUBE_LUT_BE3E 16'hBB53
`define CUBE_LUT_BE3F 16'hBB53
`define CUBE_LUT_BE40 16'hBB54
`define CUBE_LUT_BE41 16'hBB54
`define CUBE_LUT_BE42 16'hBB54
`define CUBE_LUT_BE43 16'hBB55
`define CUBE_LUT_BE44 16'hBB55
`define CUBE_LUT_BE45 16'hBB55
`define CUBE_LUT_BE46 16'hBB56
`define CUBE_LUT_BE47 16'hBB56
`define CUBE_LUT_BE48 16'hBB56
`define CUBE_LUT_BE49 16'hBB56
`define CUBE_LUT_BE4A 16'hBB57
`define CUBE_LUT_BE4B 16'hBB57
`define CUBE_LUT_BE4C 16'hBB57
`define CUBE_LUT_BE4D 16'hBB58
`define CUBE_LUT_BE4E 16'hBB58
`define CUBE_LUT_BE4F 16'hBB58
`define CUBE_LUT_BE50 16'hBB59
`define CUBE_LUT_BE51 16'hBB59
`define CUBE_LUT_BE52 16'hBB59
`define CUBE_LUT_BE53 16'hBB5A
`define CUBE_LUT_BE54 16'hBB5A
`define CUBE_LUT_BE55 16'hBB5A
`define CUBE_LUT_BE56 16'hBB5B
`define CUBE_LUT_BE57 16'hBB5B
`define CUBE_LUT_BE58 16'hBB5B
`define CUBE_LUT_BE59 16'hBB5B
`define CUBE_LUT_BE5A 16'hBB5C
`define CUBE_LUT_BE5B 16'hBB5C
`define CUBE_LUT_BE5C 16'hBB5C
`define CUBE_LUT_BE5D 16'hBB5D
`define CUBE_LUT_BE5E 16'hBB5D
`define CUBE_LUT_BE5F 16'hBB5D
`define CUBE_LUT_BE60 16'hBB5E
`define CUBE_LUT_BE61 16'hBB5E
`define CUBE_LUT_BE62 16'hBB5E
`define CUBE_LUT_BE63 16'hBB5F
`define CUBE_LUT_BE64 16'hBB5F
`define CUBE_LUT_BE65 16'hBB5F
`define CUBE_LUT_BE66 16'hBB5F
`define CUBE_LUT_BE67 16'hBB60
`define CUBE_LUT_BE68 16'hBB60
`define CUBE_LUT_BE69 16'hBB60
`define CUBE_LUT_BE6A 16'hBB61
`define CUBE_LUT_BE6B 16'hBB61
`define CUBE_LUT_BE6C 16'hBB61
`define CUBE_LUT_BE6D 16'hBB62
`define CUBE_LUT_BE6E 16'hBB62
`define CUBE_LUT_BE6F 16'hBB62
`define CUBE_LUT_BE70 16'hBB62
`define CUBE_LUT_BE71 16'hBB63
`define CUBE_LUT_BE72 16'hBB63
`define CUBE_LUT_BE73 16'hBB63
`define CUBE_LUT_BE74 16'hBB64
`define CUBE_LUT_BE75 16'hBB64
`define CUBE_LUT_BE76 16'hBB64
`define CUBE_LUT_BE77 16'hBB65
`define CUBE_LUT_BE78 16'hBB65
`define CUBE_LUT_BE79 16'hBB65
`define CUBE_LUT_BE7A 16'hBB65
`define CUBE_LUT_BE7B 16'hBB66
`define CUBE_LUT_BE7C 16'hBB66
`define CUBE_LUT_BE7D 16'hBB66
`define CUBE_LUT_BE7E 16'hBB67
`define CUBE_LUT_BE7F 16'hBB67
`define CUBE_LUT_BE80 16'hBB67
`define CUBE_LUT_BE81 16'hBB67
`define CUBE_LUT_BE82 16'hBB68
`define CUBE_LUT_BE83 16'hBB68
`define CUBE_LUT_BE84 16'hBB68
`define CUBE_LUT_BE85 16'hBB69
`define CUBE_LUT_BE86 16'hBB69
`define CUBE_LUT_BE87 16'hBB69
`define CUBE_LUT_BE88 16'hBB69
`define CUBE_LUT_BE89 16'hBB6A
`define CUBE_LUT_BE8A 16'hBB6A
`define CUBE_LUT_BE8B 16'hBB6A
`define CUBE_LUT_BE8C 16'hBB6B
`define CUBE_LUT_BE8D 16'hBB6B
`define CUBE_LUT_BE8E 16'hBB6B
`define CUBE_LUT_BE8F 16'hBB6B
`define CUBE_LUT_BE90 16'hBB6C
`define CUBE_LUT_BE91 16'hBB6C
`define CUBE_LUT_BE92 16'hBB6C
`define CUBE_LUT_BE93 16'hBB6C
`define CUBE_LUT_BE94 16'hBB6D
`define CUBE_LUT_BE95 16'hBB6D
`define CUBE_LUT_BE96 16'hBB6D
`define CUBE_LUT_BE97 16'hBB6E
`define CUBE_LUT_BE98 16'hBB6E
`define CUBE_LUT_BE99 16'hBB6E
`define CUBE_LUT_BE9A 16'hBB6E
`define CUBE_LUT_BE9B 16'hBB6F
`define CUBE_LUT_BE9C 16'hBB6F
`define CUBE_LUT_BE9D 16'hBB6F
`define CUBE_LUT_BE9E 16'hBB70
`define CUBE_LUT_BE9F 16'hBB70
`define CUBE_LUT_BEA0 16'hBB70
`define CUBE_LUT_BEA1 16'hBB70
`define CUBE_LUT_BEA2 16'hBB71
`define CUBE_LUT_BEA3 16'hBB71
`define CUBE_LUT_BEA4 16'hBB71
`define CUBE_LUT_BEA5 16'hBB71
`define CUBE_LUT_BEA6 16'hBB72
`define CUBE_LUT_BEA7 16'hBB72
`define CUBE_LUT_BEA8 16'hBB72
`define CUBE_LUT_BEA9 16'hBB72
`define CUBE_LUT_BEAA 16'hBB73
`define CUBE_LUT_BEAB 16'hBB73
`define CUBE_LUT_BEAC 16'hBB73
`define CUBE_LUT_BEAD 16'hBB74
`define CUBE_LUT_BEAE 16'hBB74
`define CUBE_LUT_BEAF 16'hBB74
`define CUBE_LUT_BEB0 16'hBB74
`define CUBE_LUT_BEB1 16'hBB75
`define CUBE_LUT_BEB2 16'hBB75
`define CUBE_LUT_BEB3 16'hBB75
`define CUBE_LUT_BEB4 16'hBB75
`define CUBE_LUT_BEB5 16'hBB76
`define CUBE_LUT_BEB6 16'hBB76
`define CUBE_LUT_BEB7 16'hBB76
`define CUBE_LUT_BEB8 16'hBB76
`define CUBE_LUT_BEB9 16'hBB77
`define CUBE_LUT_BEBA 16'hBB77
`define CUBE_LUT_BEBB 16'hBB77
`define CUBE_LUT_BEBC 16'hBB77
`define CUBE_LUT_BEBD 16'hBB78
`define CUBE_LUT_BEBE 16'hBB78
`define CUBE_LUT_BEBF 16'hBB78
`define CUBE_LUT_BEC0 16'hBB78
`define CUBE_LUT_BEC1 16'hBB79
`define CUBE_LUT_BEC2 16'hBB79
`define CUBE_LUT_BEC3 16'hBB79
`define CUBE_LUT_BEC4 16'hBB79
`define CUBE_LUT_BEC5 16'hBB7A
`define CUBE_LUT_BEC6 16'hBB7A
`define CUBE_LUT_BEC7 16'hBB7A
`define CUBE_LUT_BEC8 16'hBB7B
`define CUBE_LUT_BEC9 16'hBB7B
`define CUBE_LUT_BECA 16'hBB7B
`define CUBE_LUT_BECB 16'hBB7B
`define CUBE_LUT_BECC 16'hBB7C
`define CUBE_LUT_BECD 16'hBB7C
`define CUBE_LUT_BECE 16'hBB7C
`define CUBE_LUT_BECF 16'hBB7C
`define CUBE_LUT_BED0 16'hBB7D
`define CUBE_LUT_BED1 16'hBB7D
`define CUBE_LUT_BED2 16'hBB7D
`define CUBE_LUT_BED3 16'hBB7D
`define CUBE_LUT_BED4 16'hBB7E
`define CUBE_LUT_BED5 16'hBB7E
`define CUBE_LUT_BED6 16'hBB7E
`define CUBE_LUT_BED7 16'hBB7E
`define CUBE_LUT_BED8 16'hBB7E
`define CUBE_LUT_BED9 16'hBB7F
`define CUBE_LUT_BEDA 16'hBB7F
`define CUBE_LUT_BEDB 16'hBB7F
`define CUBE_LUT_BEDC 16'hBB7F
`define CUBE_LUT_BEDD 16'hBB80
`define CUBE_LUT_BEDE 16'hBB80
`define CUBE_LUT_BEDF 16'hBB80
`define CUBE_LUT_BEE0 16'hBB80
`define CUBE_LUT_BEE1 16'hBB81
`define CUBE_LUT_BEE2 16'hBB81
`define CUBE_LUT_BEE3 16'hBB81
`define CUBE_LUT_BEE4 16'hBB81
`define CUBE_LUT_BEE5 16'hBB82
`define CUBE_LUT_BEE6 16'hBB82
`define CUBE_LUT_BEE7 16'hBB82
`define CUBE_LUT_BEE8 16'hBB82
`define CUBE_LUT_BEE9 16'hBB83
`define CUBE_LUT_BEEA 16'hBB83
`define CUBE_LUT_BEEB 16'hBB83
`define CUBE_LUT_BEEC 16'hBB83
`define CUBE_LUT_BEED 16'hBB84
`define CUBE_LUT_BEEE 16'hBB84
`define CUBE_LUT_BEEF 16'hBB84
`define CUBE_LUT_BEF0 16'hBB84
`define CUBE_LUT_BEF1 16'hBB84
`define CUBE_LUT_BEF2 16'hBB85
`define CUBE_LUT_BEF3 16'hBB85
`define CUBE_LUT_BEF4 16'hBB85
`define CUBE_LUT_BEF5 16'hBB85
`define CUBE_LUT_BEF6 16'hBB86
`define CUBE_LUT_BEF7 16'hBB86
`define CUBE_LUT_BEF8 16'hBB86
`define CUBE_LUT_BEF9 16'hBB86
`define CUBE_LUT_BEFA 16'hBB87
`define CUBE_LUT_BEFB 16'hBB87
`define CUBE_LUT_BEFC 16'hBB87
`define CUBE_LUT_BEFD 16'hBB87
`define CUBE_LUT_BEFE 16'hBB87
`define CUBE_LUT_BEFF 16'hBB88
`define CUBE_LUT_BF00 16'hBB88
`define CUBE_LUT_BF01 16'hBB88
`define CUBE_LUT_BF02 16'hBB88
`define CUBE_LUT_BF03 16'hBB89
`define CUBE_LUT_BF04 16'hBB89
`define CUBE_LUT_BF05 16'hBB89
`define CUBE_LUT_BF06 16'hBB89
`define CUBE_LUT_BF07 16'hBB8A
`define CUBE_LUT_BF08 16'hBB8A
`define CUBE_LUT_BF09 16'hBB8A
`define CUBE_LUT_BF0A 16'hBB8A
`define CUBE_LUT_BF0B 16'hBB8A
`define CUBE_LUT_BF0C 16'hBB8B
`define CUBE_LUT_BF0D 16'hBB8B
`define CUBE_LUT_BF0E 16'hBB8B
`define CUBE_LUT_BF0F 16'hBB8B
`define CUBE_LUT_BF10 16'hBB8C
`define CUBE_LUT_BF11 16'hBB8C
`define CUBE_LUT_BF12 16'hBB8C
`define CUBE_LUT_BF13 16'hBB8C
`define CUBE_LUT_BF14 16'hBB8C
`define CUBE_LUT_BF15 16'hBB8D
`define CUBE_LUT_BF16 16'hBB8D
`define CUBE_LUT_BF17 16'hBB8D
`define CUBE_LUT_BF18 16'hBB8D
`define CUBE_LUT_BF19 16'hBB8D
`define CUBE_LUT_BF1A 16'hBB8E
`define CUBE_LUT_BF1B 16'hBB8E
`define CUBE_LUT_BF1C 16'hBB8E
`define CUBE_LUT_BF1D 16'hBB8E
`define CUBE_LUT_BF1E 16'hBB8F
`define CUBE_LUT_BF1F 16'hBB8F
`define CUBE_LUT_BF20 16'hBB8F
`define CUBE_LUT_BF21 16'hBB8F
`define CUBE_LUT_BF22 16'hBB8F
`define CUBE_LUT_BF23 16'hBB90
`define CUBE_LUT_BF24 16'hBB90
`define CUBE_LUT_BF25 16'hBB90
`define CUBE_LUT_BF26 16'hBB90
`define CUBE_LUT_BF27 16'hBB91
`define CUBE_LUT_BF28 16'hBB91
`define CUBE_LUT_BF29 16'hBB91
`define CUBE_LUT_BF2A 16'hBB91
`define CUBE_LUT_BF2B 16'hBB91
`define CUBE_LUT_BF2C 16'hBB92
`define CUBE_LUT_BF2D 16'hBB92
`define CUBE_LUT_BF2E 16'hBB92
`define CUBE_LUT_BF2F 16'hBB92
`define CUBE_LUT_BF30 16'hBB92
`define CUBE_LUT_BF31 16'hBB93
`define CUBE_LUT_BF32 16'hBB93
`define CUBE_LUT_BF33 16'hBB93
`define CUBE_LUT_BF34 16'hBB93
`define CUBE_LUT_BF35 16'hBB93
`define CUBE_LUT_BF36 16'hBB94
`define CUBE_LUT_BF37 16'hBB94
`define CUBE_LUT_BF38 16'hBB94
`define CUBE_LUT_BF39 16'hBB94
`define CUBE_LUT_BF3A 16'hBB94
`define CUBE_LUT_BF3B 16'hBB95
`define CUBE_LUT_BF3C 16'hBB95
`define CUBE_LUT_BF3D 16'hBB95
`define CUBE_LUT_BF3E 16'hBB95
`define CUBE_LUT_BF3F 16'hBB95
`define CUBE_LUT_BF40 16'hBB96
`define CUBE_LUT_BF41 16'hBB96
`define CUBE_LUT_BF42 16'hBB96
`define CUBE_LUT_BF43 16'hBB96
`define CUBE_LUT_BF44 16'hBB96
`define CUBE_LUT_BF45 16'hBB97
`define CUBE_LUT_BF46 16'hBB97
`define CUBE_LUT_BF47 16'hBB97
`define CUBE_LUT_BF48 16'hBB97
`define CUBE_LUT_BF49 16'hBB97
`define CUBE_LUT_BF4A 16'hBB98
`define CUBE_LUT_BF4B 16'hBB98
`define CUBE_LUT_BF4C 16'hBB98
`define CUBE_LUT_BF4D 16'hBB98
`define CUBE_LUT_BF4E 16'hBB98
`define CUBE_LUT_BF4F 16'hBB99
`define CUBE_LUT_BF50 16'hBB99
`define CUBE_LUT_BF51 16'hBB99
`define CUBE_LUT_BF52 16'hBB99
`define CUBE_LUT_BF53 16'hBB99
`define CUBE_LUT_BF54 16'hBB9A
`define CUBE_LUT_BF55 16'hBB9A
`define CUBE_LUT_BF56 16'hBB9A
`define CUBE_LUT_BF57 16'hBB9A
`define CUBE_LUT_BF58 16'hBB9A
`define CUBE_LUT_BF59 16'hBB9B
`define CUBE_LUT_BF5A 16'hBB9B
`define CUBE_LUT_BF5B 16'hBB9B
`define CUBE_LUT_BF5C 16'hBB9B
`define CUBE_LUT_BF5D 16'hBB9B
`define CUBE_LUT_BF5E 16'hBB9C
`define CUBE_LUT_BF5F 16'hBB9C
`define CUBE_LUT_BF60 16'hBB9C
`define CUBE_LUT_BF61 16'hBB9C
`define CUBE_LUT_BF62 16'hBB9C
`define CUBE_LUT_BF63 16'hBB9D
`define CUBE_LUT_BF64 16'hBB9D
`define CUBE_LUT_BF65 16'hBB9D
`define CUBE_LUT_BF66 16'hBB9D
`define CUBE_LUT_BF67 16'hBB9D
`define CUBE_LUT_BF68 16'hBB9D
`define CUBE_LUT_BF69 16'hBB9E
`define CUBE_LUT_BF6A 16'hBB9E
`define CUBE_LUT_BF6B 16'hBB9E
`define CUBE_LUT_BF6C 16'hBB9E
`define CUBE_LUT_BF6D 16'hBB9E
`define CUBE_LUT_BF6E 16'hBB9F
`define CUBE_LUT_BF6F 16'hBB9F
`define CUBE_LUT_BF70 16'hBB9F
`define CUBE_LUT_BF71 16'hBB9F
`define CUBE_LUT_BF72 16'hBB9F
`define CUBE_LUT_BF73 16'hBBA0
`define CUBE_LUT_BF74 16'hBBA0
`define CUBE_LUT_BF75 16'hBBA0
`define CUBE_LUT_BF76 16'hBBA0
`define CUBE_LUT_BF77 16'hBBA0
`define CUBE_LUT_BF78 16'hBBA0
`define CUBE_LUT_BF79 16'hBBA1
`define CUBE_LUT_BF7A 16'hBBA1
`define CUBE_LUT_BF7B 16'hBBA1
`define CUBE_LUT_BF7C 16'hBBA1
`define CUBE_LUT_BF7D 16'hBBA1
`define CUBE_LUT_BF7E 16'hBBA2
`define CUBE_LUT_BF7F 16'hBBA2
`define CUBE_LUT_BF80 16'hBBA2
`define CUBE_LUT_BF81 16'hBBA2
`define CUBE_LUT_BF82 16'hBBA2
`define CUBE_LUT_BF83 16'hBBA2
`define CUBE_LUT_BF84 16'hBBA3
`define CUBE_LUT_BF85 16'hBBA3
`define CUBE_LUT_BF86 16'hBBA3
`define CUBE_LUT_BF87 16'hBBA3
`define CUBE_LUT_BF88 16'hBBA3
`define CUBE_LUT_BF89 16'hBBA3
`define CUBE_LUT_BF8A 16'hBBA4
`define CUBE_LUT_BF8B 16'hBBA4
`define CUBE_LUT_BF8C 16'hBBA4
`define CUBE_LUT_BF8D 16'hBBA4
`define CUBE_LUT_BF8E 16'hBBA4
`define CUBE_LUT_BF8F 16'hBBA5
`define CUBE_LUT_BF90 16'hBBA5
`define CUBE_LUT_BF91 16'hBBA5
`define CUBE_LUT_BF92 16'hBBA5
`define CUBE_LUT_BF93 16'hBBA5
`define CUBE_LUT_BF94 16'hBBA5
`define CUBE_LUT_BF95 16'hBBA6
`define CUBE_LUT_BF96 16'hBBA6
`define CUBE_LUT_BF97 16'hBBA6
`define CUBE_LUT_BF98 16'hBBA6
`define CUBE_LUT_BF99 16'hBBA6
`define CUBE_LUT_BF9A 16'hBBA6
`define CUBE_LUT_BF9B 16'hBBA7
`define CUBE_LUT_BF9C 16'hBBA7
`define CUBE_LUT_BF9D 16'hBBA7
`define CUBE_LUT_BF9E 16'hBBA7
`define CUBE_LUT_BF9F 16'hBBA7
`define CUBE_LUT_BFA0 16'hBBA7
`define CUBE_LUT_BFA1 16'hBBA8
`define CUBE_LUT_BFA2 16'hBBA8
`define CUBE_LUT_BFA3 16'hBBA8
`define CUBE_LUT_BFA4 16'hBBA8
`define CUBE_LUT_BFA5 16'hBBA8
`define CUBE_LUT_BFA6 16'hBBA8
`define CUBE_LUT_BFA7 16'hBBA9
`define CUBE_LUT_BFA8 16'hBBA9
`define CUBE_LUT_BFA9 16'hBBA9
`define CUBE_LUT_BFAA 16'hBBA9
`define CUBE_LUT_BFAB 16'hBBA9
`define CUBE_LUT_BFAC 16'hBBA9
`define CUBE_LUT_BFAD 16'hBBAA
`define CUBE_LUT_BFAE 16'hBBAA
`define CUBE_LUT_BFAF 16'hBBAA
`define CUBE_LUT_BFB0 16'hBBAA
`define CUBE_LUT_BFB1 16'hBBAA
`define CUBE_LUT_BFB2 16'hBBAA
`define CUBE_LUT_BFB3 16'hBBAB
`define CUBE_LUT_BFB4 16'hBBAB
`define CUBE_LUT_BFB5 16'hBBAB
`define CUBE_LUT_BFB6 16'hBBAB
`define CUBE_LUT_BFB7 16'hBBAB
`define CUBE_LUT_BFB8 16'hBBAB
`define CUBE_LUT_BFB9 16'hBBAC
`define CUBE_LUT_BFBA 16'hBBAC
`define CUBE_LUT_BFBB 16'hBBAC
`define CUBE_LUT_BFBC 16'hBBAC
`define CUBE_LUT_BFBD 16'hBBAC
`define CUBE_LUT_BFBE 16'hBBAC
`define CUBE_LUT_BFBF 16'hBBAD
`define CUBE_LUT_BFC0 16'hBBAD
`define CUBE_LUT_BFC1 16'hBBAD
`define CUBE_LUT_BFC2 16'hBBAD
`define CUBE_LUT_BFC3 16'hBBAD
`define CUBE_LUT_BFC4 16'hBBAD
`define CUBE_LUT_BFC5 16'hBBAE
`define CUBE_LUT_BFC6 16'hBBAE
`define CUBE_LUT_BFC7 16'hBBAE
`define CUBE_LUT_BFC8 16'hBBAE
`define CUBE_LUT_BFC9 16'hBBAE
`define CUBE_LUT_BFCA 16'hBBAE
`define CUBE_LUT_BFCB 16'hBBAE
`define CUBE_LUT_BFCC 16'hBBAF
`define CUBE_LUT_BFCD 16'hBBAF
`define CUBE_LUT_BFCE 16'hBBAF
`define CUBE_LUT_BFCF 16'hBBAF
`define CUBE_LUT_BFD0 16'hBBAF
`define CUBE_LUT_BFD1 16'hBBAF
`define CUBE_LUT_BFD2 16'hBBB0
`define CUBE_LUT_BFD3 16'hBBB0
`define CUBE_LUT_BFD4 16'hBBB0
`define CUBE_LUT_BFD5 16'hBBB0
`define CUBE_LUT_BFD6 16'hBBB0
`define CUBE_LUT_BFD7 16'hBBB0
`define CUBE_LUT_BFD8 16'hBBB0
`define CUBE_LUT_BFD9 16'hBBB1
`define CUBE_LUT_BFDA 16'hBBB1
`define CUBE_LUT_BFDB 16'hBBB1
`define CUBE_LUT_BFDC 16'hBBB1
`define CUBE_LUT_BFDD 16'hBBB1
`define CUBE_LUT_BFDE 16'hBBB1
`define CUBE_LUT_BFDF 16'hBBB2
`define CUBE_LUT_BFE0 16'hBBB2
`define CUBE_LUT_BFE1 16'hBBB2
`define CUBE_LUT_BFE2 16'hBBB2
`define CUBE_LUT_BFE3 16'hBBB2
`define CUBE_LUT_BFE4 16'hBBB2
`define CUBE_LUT_BFE5 16'hBBB2
`define CUBE_LUT_BFE6 16'hBBB3
`define CUBE_LUT_BFE7 16'hBBB3
`define CUBE_LUT_BFE8 16'hBBB3
`define CUBE_LUT_BFE9 16'hBBB3
`define CUBE_LUT_BFEA 16'hBBB3
`define CUBE_LUT_BFEB 16'hBBB3
`define CUBE_LUT_BFEC 16'hBBB3
`define CUBE_LUT_BFED 16'hBBB4
`define CUBE_LUT_BFEE 16'hBBB4
`define CUBE_LUT_BFEF 16'hBBB4
`define CUBE_LUT_BFF0 16'hBBB4
`define CUBE_LUT_BFF1 16'hBBB4
`define CUBE_LUT_BFF2 16'hBBB4
`define CUBE_LUT_BFF3 16'hBBB4
`define CUBE_LUT_BFF4 16'hBBB5
`define CUBE_LUT_BFF5 16'hBBB5
`define CUBE_LUT_BFF6 16'hBBB5
`define CUBE_LUT_BFF7 16'hBBB5
`define CUBE_LUT_BFF8 16'hBBB5
`define CUBE_LUT_BFF9 16'hBBB5
`define CUBE_LUT_BFFA 16'hBBB5
`define CUBE_LUT_BFFB 16'hBBB6
`define CUBE_LUT_BFFC 16'hBBB6
`define CUBE_LUT_BFFD 16'hBBB6
`define CUBE_LUT_BFFE 16'hBBB6
`define CUBE_LUT_BFFF 16'hBBB6
`define CUBE_LUT_C000 16'hBBB6
`define CUBE_LUT_C001 16'hBBB7
`define CUBE_LUT_C002 16'hBBB7
`define CUBE_LUT_C003 16'hBBB7
`define CUBE_LUT_C004 16'hBBB7
`define CUBE_LUT_C005 16'hBBB8
`define CUBE_LUT_C006 16'hBBB8
`define CUBE_LUT_C007 16'hBBB8
`define CUBE_LUT_C008 16'hBBB9
`define CUBE_LUT_C009 16'hBBB9
`define CUBE_LUT_C00A 16'hBBB9
`define CUBE_LUT_C00B 16'hBBB9
`define CUBE_LUT_C00C 16'hBBBA
`define CUBE_LUT_C00D 16'hBBBA
`define CUBE_LUT_C00E 16'hBBBA
`define CUBE_LUT_C00F 16'hBBBA
`define CUBE_LUT_C010 16'hBBBB
`define CUBE_LUT_C011 16'hBBBB
`define CUBE_LUT_C012 16'hBBBB
`define CUBE_LUT_C013 16'hBBBC
`define CUBE_LUT_C014 16'hBBBC
`define CUBE_LUT_C015 16'hBBBC
`define CUBE_LUT_C016 16'hBBBC
`define CUBE_LUT_C017 16'hBBBD
`define CUBE_LUT_C018 16'hBBBD
`define CUBE_LUT_C019 16'hBBBD
`define CUBE_LUT_C01A 16'hBBBD
`define CUBE_LUT_C01B 16'hBBBE
`define CUBE_LUT_C01C 16'hBBBE
`define CUBE_LUT_C01D 16'hBBBE
`define CUBE_LUT_C01E 16'hBBBE
`define CUBE_LUT_C01F 16'hBBBF
`define CUBE_LUT_C020 16'hBBBF
`define CUBE_LUT_C021 16'hBBBF
`define CUBE_LUT_C022 16'hBBBF
`define CUBE_LUT_C023 16'hBBC0
`define CUBE_LUT_C024 16'hBBC0
`define CUBE_LUT_C025 16'hBBC0
`define CUBE_LUT_C026 16'hBBC0
`define CUBE_LUT_C027 16'hBBC1
`define CUBE_LUT_C028 16'hBBC1
`define CUBE_LUT_C029 16'hBBC1
`define CUBE_LUT_C02A 16'hBBC1
`define CUBE_LUT_C02B 16'hBBC2
`define CUBE_LUT_C02C 16'hBBC2
`define CUBE_LUT_C02D 16'hBBC2
`define CUBE_LUT_C02E 16'hBBC2
`define CUBE_LUT_C02F 16'hBBC2
`define CUBE_LUT_C030 16'hBBC3
`define CUBE_LUT_C031 16'hBBC3
`define CUBE_LUT_C032 16'hBBC3
`define CUBE_LUT_C033 16'hBBC3
`define CUBE_LUT_C034 16'hBBC4
`define CUBE_LUT_C035 16'hBBC4
`define CUBE_LUT_C036 16'hBBC4
`define CUBE_LUT_C037 16'hBBC4
`define CUBE_LUT_C038 16'hBBC5
`define CUBE_LUT_C039 16'hBBC5
`define CUBE_LUT_C03A 16'hBBC5
`define CUBE_LUT_C03B 16'hBBC5
`define CUBE_LUT_C03C 16'hBBC6
`define CUBE_LUT_C03D 16'hBBC6
`define CUBE_LUT_C03E 16'hBBC6
`define CUBE_LUT_C03F 16'hBBC6
`define CUBE_LUT_C040 16'hBBC6
`define CUBE_LUT_C041 16'hBBC7
`define CUBE_LUT_C042 16'hBBC7
`define CUBE_LUT_C043 16'hBBC7
`define CUBE_LUT_C044 16'hBBC7
`define CUBE_LUT_C045 16'hBBC7
`define CUBE_LUT_C046 16'hBBC8
`define CUBE_LUT_C047 16'hBBC8
`define CUBE_LUT_C048 16'hBBC8
`define CUBE_LUT_C049 16'hBBC8
`define CUBE_LUT_C04A 16'hBBC9
`define CUBE_LUT_C04B 16'hBBC9
`define CUBE_LUT_C04C 16'hBBC9
`define CUBE_LUT_C04D 16'hBBC9
`define CUBE_LUT_C04E 16'hBBC9
`define CUBE_LUT_C04F 16'hBBCA
`define CUBE_LUT_C050 16'hBBCA
`define CUBE_LUT_C051 16'hBBCA
`define CUBE_LUT_C052 16'hBBCA
`define CUBE_LUT_C053 16'hBBCA
`define CUBE_LUT_C054 16'hBBCB
`define CUBE_LUT_C055 16'hBBCB
`define CUBE_LUT_C056 16'hBBCB
`define CUBE_LUT_C057 16'hBBCB
`define CUBE_LUT_C058 16'hBBCB
`define CUBE_LUT_C059 16'hBBCC
`define CUBE_LUT_C05A 16'hBBCC
`define CUBE_LUT_C05B 16'hBBCC
`define CUBE_LUT_C05C 16'hBBCC
`define CUBE_LUT_C05D 16'hBBCC
`define CUBE_LUT_C05E 16'hBBCD
`define CUBE_LUT_C05F 16'hBBCD
`define CUBE_LUT_C060 16'hBBCD
`define CUBE_LUT_C061 16'hBBCD
`define CUBE_LUT_C062 16'hBBCD
`define CUBE_LUT_C063 16'hBBCE
`define CUBE_LUT_C064 16'hBBCE
`define CUBE_LUT_C065 16'hBBCE
`define CUBE_LUT_C066 16'hBBCE
`define CUBE_LUT_C067 16'hBBCE
`define CUBE_LUT_C068 16'hBBCF
`define CUBE_LUT_C069 16'hBBCF
`define CUBE_LUT_C06A 16'hBBCF
`define CUBE_LUT_C06B 16'hBBCF
`define CUBE_LUT_C06C 16'hBBCF
`define CUBE_LUT_C06D 16'hBBD0
`define CUBE_LUT_C06E 16'hBBD0
`define CUBE_LUT_C06F 16'hBBD0
`define CUBE_LUT_C070 16'hBBD0
`define CUBE_LUT_C071 16'hBBD0
`define CUBE_LUT_C072 16'hBBD0
`define CUBE_LUT_C073 16'hBBD1
`define CUBE_LUT_C074 16'hBBD1
`define CUBE_LUT_C075 16'hBBD1
`define CUBE_LUT_C076 16'hBBD1
`define CUBE_LUT_C077 16'hBBD1
`define CUBE_LUT_C078 16'hBBD2
`define CUBE_LUT_C079 16'hBBD2
`define CUBE_LUT_C07A 16'hBBD2
`define CUBE_LUT_C07B 16'hBBD2
`define CUBE_LUT_C07C 16'hBBD2
`define CUBE_LUT_C07D 16'hBBD2
`define CUBE_LUT_C07E 16'hBBD3
`define CUBE_LUT_C07F 16'hBBD3
`define CUBE_LUT_C080 16'hBBD3
`define CUBE_LUT_C081 16'hBBD3
`define CUBE_LUT_C082 16'hBBD3
`define CUBE_LUT_C083 16'hBBD4
`define CUBE_LUT_C084 16'hBBD4
`define CUBE_LUT_C085 16'hBBD4
`define CUBE_LUT_C086 16'hBBD4
`define CUBE_LUT_C087 16'hBBD4
`define CUBE_LUT_C088 16'hBBD4
`define CUBE_LUT_C089 16'hBBD5
`define CUBE_LUT_C08A 16'hBBD5
`define CUBE_LUT_C08B 16'hBBD5
`define CUBE_LUT_C08C 16'hBBD5
`define CUBE_LUT_C08D 16'hBBD5
`define CUBE_LUT_C08E 16'hBBD5
`define CUBE_LUT_C08F 16'hBBD6
`define CUBE_LUT_C090 16'hBBD6
`define CUBE_LUT_C091 16'hBBD6
`define CUBE_LUT_C092 16'hBBD6
`define CUBE_LUT_C093 16'hBBD6
`define CUBE_LUT_C094 16'hBBD6
`define CUBE_LUT_C095 16'hBBD7
`define CUBE_LUT_C096 16'hBBD7
`define CUBE_LUT_C097 16'hBBD7
`define CUBE_LUT_C098 16'hBBD7
`define CUBE_LUT_C099 16'hBBD7
`define CUBE_LUT_C09A 16'hBBD7
`define CUBE_LUT_C09B 16'hBBD7
`define CUBE_LUT_C09C 16'hBBD8
`define CUBE_LUT_C09D 16'hBBD8
`define CUBE_LUT_C09E 16'hBBD8
`define CUBE_LUT_C09F 16'hBBD8
`define CUBE_LUT_C0A0 16'hBBD8
`define CUBE_LUT_C0A1 16'hBBD8
`define CUBE_LUT_C0A2 16'hBBD9
`define CUBE_LUT_C0A3 16'hBBD9
`define CUBE_LUT_C0A4 16'hBBD9
`define CUBE_LUT_C0A5 16'hBBD9
`define CUBE_LUT_C0A6 16'hBBD9
`define CUBE_LUT_C0A7 16'hBBD9
`define CUBE_LUT_C0A8 16'hBBD9
`define CUBE_LUT_C0A9 16'hBBDA
`define CUBE_LUT_C0AA 16'hBBDA
`define CUBE_LUT_C0AB 16'hBBDA
`define CUBE_LUT_C0AC 16'hBBDA
`define CUBE_LUT_C0AD 16'hBBDA
`define CUBE_LUT_C0AE 16'hBBDA
`define CUBE_LUT_C0AF 16'hBBDA
`define CUBE_LUT_C0B0 16'hBBDB
`define CUBE_LUT_C0B1 16'hBBDB
`define CUBE_LUT_C0B2 16'hBBDB
`define CUBE_LUT_C0B3 16'hBBDB
`define CUBE_LUT_C0B4 16'hBBDB
`define CUBE_LUT_C0B5 16'hBBDB
`define CUBE_LUT_C0B6 16'hBBDB
`define CUBE_LUT_C0B7 16'hBBDC
`define CUBE_LUT_C0B8 16'hBBDC
`define CUBE_LUT_C0B9 16'hBBDC
`define CUBE_LUT_C0BA 16'hBBDC
`define CUBE_LUT_C0BB 16'hBBDC
`define CUBE_LUT_C0BC 16'hBBDC
`define CUBE_LUT_C0BD 16'hBBDC
`define CUBE_LUT_C0BE 16'hBBDD
`define CUBE_LUT_C0BF 16'hBBDD
`define CUBE_LUT_C0C0 16'hBBDD
`define CUBE_LUT_C0C1 16'hBBDD
`define CUBE_LUT_C0C2 16'hBBDD
`define CUBE_LUT_C0C3 16'hBBDD
`define CUBE_LUT_C0C4 16'hBBDD
`define CUBE_LUT_C0C5 16'hBBDE
`define CUBE_LUT_C0C6 16'hBBDE
`define CUBE_LUT_C0C7 16'hBBDE
`define CUBE_LUT_C0C8 16'hBBDE
`define CUBE_LUT_C0C9 16'hBBDE
`define CUBE_LUT_C0CA 16'hBBDE
`define CUBE_LUT_C0CB 16'hBBDE
`define CUBE_LUT_C0CC 16'hBBDE
`define CUBE_LUT_C0CD 16'hBBDF
`define CUBE_LUT_C0CE 16'hBBDF
`define CUBE_LUT_C0CF 16'hBBDF
`define CUBE_LUT_C0D0 16'hBBDF
`define CUBE_LUT_C0D1 16'hBBDF
`define CUBE_LUT_C0D2 16'hBBDF
`define CUBE_LUT_C0D3 16'hBBDF
`define CUBE_LUT_C0D4 16'hBBDF
`define CUBE_LUT_C0D5 16'hBBE0
`define CUBE_LUT_C0D6 16'hBBE0
`define CUBE_LUT_C0D7 16'hBBE0
`define CUBE_LUT_C0D8 16'hBBE0
`define CUBE_LUT_C0D9 16'hBBE0
`define CUBE_LUT_C0DA 16'hBBE0
`define CUBE_LUT_C0DB 16'hBBE0
`define CUBE_LUT_C0DC 16'hBBE0
`define CUBE_LUT_C0DD 16'hBBE1
`define CUBE_LUT_C0DE 16'hBBE1
`define CUBE_LUT_C0DF 16'hBBE1
`define CUBE_LUT_C0E0 16'hBBE1
`define CUBE_LUT_C0E1 16'hBBE1
`define CUBE_LUT_C0E2 16'hBBE1
`define CUBE_LUT_C0E3 16'hBBE1
`define CUBE_LUT_C0E4 16'hBBE1
`define CUBE_LUT_C0E5 16'hBBE2
`define CUBE_LUT_C0E6 16'hBBE2
`define CUBE_LUT_C0E7 16'hBBE2
`define CUBE_LUT_C0E8 16'hBBE2
`define CUBE_LUT_C0E9 16'hBBE2
`define CUBE_LUT_C0EA 16'hBBE2
`define CUBE_LUT_C0EB 16'hBBE2
`define CUBE_LUT_C0EC 16'hBBE2
`define CUBE_LUT_C0ED 16'hBBE2
`define CUBE_LUT_C0EE 16'hBBE3
`define CUBE_LUT_C0EF 16'hBBE3
`define CUBE_LUT_C0F0 16'hBBE3
`define CUBE_LUT_C0F1 16'hBBE3
`define CUBE_LUT_C0F2 16'hBBE3
`define CUBE_LUT_C0F3 16'hBBE3
`define CUBE_LUT_C0F4 16'hBBE3
`define CUBE_LUT_C0F5 16'hBBE3
`define CUBE_LUT_C0F6 16'hBBE4
`define CUBE_LUT_C0F7 16'hBBE4
`define CUBE_LUT_C0F8 16'hBBE4
`define CUBE_LUT_C0F9 16'hBBE4
`define CUBE_LUT_C0FA 16'hBBE4
`define CUBE_LUT_C0FB 16'hBBE4
`define CUBE_LUT_C0FC 16'hBBE4
`define CUBE_LUT_C0FD 16'hBBE4
`define CUBE_LUT_C0FE 16'hBBE4
`define CUBE_LUT_C0FF 16'hBBE4
`define CUBE_LUT_C100 16'hBBE5
`define CUBE_LUT_C101 16'hBBE5
`define CUBE_LUT_C102 16'hBBE5
`define CUBE_LUT_C103 16'hBBE5
`define CUBE_LUT_C104 16'hBBE5
`define CUBE_LUT_C105 16'hBBE5
`define CUBE_LUT_C106 16'hBBE5
`define CUBE_LUT_C107 16'hBBE5
`define CUBE_LUT_C108 16'hBBE5
`define CUBE_LUT_C109 16'hBBE6
`define CUBE_LUT_C10A 16'hBBE6
`define CUBE_LUT_C10B 16'hBBE6
`define CUBE_LUT_C10C 16'hBBE6
`define CUBE_LUT_C10D 16'hBBE6
`define CUBE_LUT_C10E 16'hBBE6
`define CUBE_LUT_C10F 16'hBBE6
`define CUBE_LUT_C110 16'hBBE6
`define CUBE_LUT_C111 16'hBBE6
`define CUBE_LUT_C112 16'hBBE6
`define CUBE_LUT_C113 16'hBBE7
`define CUBE_LUT_C114 16'hBBE7
`define CUBE_LUT_C115 16'hBBE7
`define CUBE_LUT_C116 16'hBBE7
`define CUBE_LUT_C117 16'hBBE7
`define CUBE_LUT_C118 16'hBBE7
`define CUBE_LUT_C119 16'hBBE7
`define CUBE_LUT_C11A 16'hBBE7
`define CUBE_LUT_C11B 16'hBBE7
`define CUBE_LUT_C11C 16'hBBE7
`define CUBE_LUT_C11D 16'hBBE8
`define CUBE_LUT_C11E 16'hBBE8
`define CUBE_LUT_C11F 16'hBBE8
`define CUBE_LUT_C120 16'hBBE8
`define CUBE_LUT_C121 16'hBBE8
`define CUBE_LUT_C122 16'hBBE8
`define CUBE_LUT_C123 16'hBBE8
`define CUBE_LUT_C124 16'hBBE8
`define CUBE_LUT_C125 16'hBBE8
`define CUBE_LUT_C126 16'hBBE8
`define CUBE_LUT_C127 16'hBBE8
`define CUBE_LUT_C128 16'hBBE9
`define CUBE_LUT_C129 16'hBBE9
`define CUBE_LUT_C12A 16'hBBE9
`define CUBE_LUT_C12B 16'hBBE9
`define CUBE_LUT_C12C 16'hBBE9
`define CUBE_LUT_C12D 16'hBBE9
`define CUBE_LUT_C12E 16'hBBE9
`define CUBE_LUT_C12F 16'hBBE9
`define CUBE_LUT_C130 16'hBBE9
`define CUBE_LUT_C131 16'hBBE9
`define CUBE_LUT_C132 16'hBBE9
`define CUBE_LUT_C133 16'hBBEA
`define CUBE_LUT_C134 16'hBBEA
`define CUBE_LUT_C135 16'hBBEA
`define CUBE_LUT_C136 16'hBBEA
`define CUBE_LUT_C137 16'hBBEA
`define CUBE_LUT_C138 16'hBBEA
`define CUBE_LUT_C139 16'hBBEA
`define CUBE_LUT_C13A 16'hBBEA
`define CUBE_LUT_C13B 16'hBBEA
`define CUBE_LUT_C13C 16'hBBEA
`define CUBE_LUT_C13D 16'hBBEA
`define CUBE_LUT_C13E 16'hBBEA
`define CUBE_LUT_C13F 16'hBBEB
`define CUBE_LUT_C140 16'hBBEB
`define CUBE_LUT_C141 16'hBBEB
`define CUBE_LUT_C142 16'hBBEB
`define CUBE_LUT_C143 16'hBBEB
`define CUBE_LUT_C144 16'hBBEB
`define CUBE_LUT_C145 16'hBBEB
`define CUBE_LUT_C146 16'hBBEB
`define CUBE_LUT_C147 16'hBBEB
`define CUBE_LUT_C148 16'hBBEB
`define CUBE_LUT_C149 16'hBBEB
`define CUBE_LUT_C14A 16'hBBEB
`define CUBE_LUT_C14B 16'hBBEC
`define CUBE_LUT_C14C 16'hBBEC
`define CUBE_LUT_C14D 16'hBBEC
`define CUBE_LUT_C14E 16'hBBEC
`define CUBE_LUT_C14F 16'hBBEC
`define CUBE_LUT_C150 16'hBBEC
`define CUBE_LUT_C151 16'hBBEC
`define CUBE_LUT_C152 16'hBBEC
`define CUBE_LUT_C153 16'hBBEC
`define CUBE_LUT_C154 16'hBBEC
`define CUBE_LUT_C155 16'hBBEC
`define CUBE_LUT_C156 16'hBBEC
`define CUBE_LUT_C157 16'hBBEC
`define CUBE_LUT_C158 16'hBBED
`define CUBE_LUT_C159 16'hBBED
`define CUBE_LUT_C15A 16'hBBED
`define CUBE_LUT_C15B 16'hBBED
`define CUBE_LUT_C15C 16'hBBED
`define CUBE_LUT_C15D 16'hBBED
`define CUBE_LUT_C15E 16'hBBED
`define CUBE_LUT_C15F 16'hBBED
`define CUBE_LUT_C160 16'hBBED
`define CUBE_LUT_C161 16'hBBED
`define CUBE_LUT_C162 16'hBBED
`define CUBE_LUT_C163 16'hBBED
`define CUBE_LUT_C164 16'hBBED
`define CUBE_LUT_C165 16'hBBED
`define CUBE_LUT_C166 16'hBBEE
`define CUBE_LUT_C167 16'hBBEE
`define CUBE_LUT_C168 16'hBBEE
`define CUBE_LUT_C169 16'hBBEE
`define CUBE_LUT_C16A 16'hBBEE
`define CUBE_LUT_C16B 16'hBBEE
`define CUBE_LUT_C16C 16'hBBEE
`define CUBE_LUT_C16D 16'hBBEE
`define CUBE_LUT_C16E 16'hBBEE
`define CUBE_LUT_C16F 16'hBBEE
`define CUBE_LUT_C170 16'hBBEE
`define CUBE_LUT_C171 16'hBBEE
`define CUBE_LUT_C172 16'hBBEE
`define CUBE_LUT_C173 16'hBBEE
`define CUBE_LUT_C174 16'hBBEF
`define CUBE_LUT_C175 16'hBBEF
`define CUBE_LUT_C176 16'hBBEF
`define CUBE_LUT_C177 16'hBBEF
`define CUBE_LUT_C178 16'hBBEF
`define CUBE_LUT_C179 16'hBBEF
`define CUBE_LUT_C17A 16'hBBEF
`define CUBE_LUT_C17B 16'hBBEF
`define CUBE_LUT_C17C 16'hBBEF
`define CUBE_LUT_C17D 16'hBBEF
`define CUBE_LUT_C17E 16'hBBEF
`define CUBE_LUT_C17F 16'hBBEF
`define CUBE_LUT_C180 16'hBBEF
`define CUBE_LUT_C181 16'hBBEF
`define CUBE_LUT_C182 16'hBBEF
`define CUBE_LUT_C183 16'hBBF0
`define CUBE_LUT_C184 16'hBBF0
`define CUBE_LUT_C185 16'hBBF0
`define CUBE_LUT_C186 16'hBBF0
`define CUBE_LUT_C187 16'hBBF0
`define CUBE_LUT_C188 16'hBBF0
`define CUBE_LUT_C189 16'hBBF0
`define CUBE_LUT_C18A 16'hBBF0
`define CUBE_LUT_C18B 16'hBBF0
`define CUBE_LUT_C18C 16'hBBF0
`define CUBE_LUT_C18D 16'hBBF0
`define CUBE_LUT_C18E 16'hBBF0
`define CUBE_LUT_C18F 16'hBBF0
`define CUBE_LUT_C190 16'hBBF0
`define CUBE_LUT_C191 16'hBBF0
`define CUBE_LUT_C192 16'hBBF0
`define CUBE_LUT_C193 16'hBBF1
`define CUBE_LUT_C194 16'hBBF1
`define CUBE_LUT_C195 16'hBBF1
`define CUBE_LUT_C196 16'hBBF1
`define CUBE_LUT_C197 16'hBBF1
`define CUBE_LUT_C198 16'hBBF1
`define CUBE_LUT_C199 16'hBBF1
`define CUBE_LUT_C19A 16'hBBF1
`define CUBE_LUT_C19B 16'hBBF1
`define CUBE_LUT_C19C 16'hBBF1
`define CUBE_LUT_C19D 16'hBBF1
`define CUBE_LUT_C19E 16'hBBF1
`define CUBE_LUT_C19F 16'hBBF1
`define CUBE_LUT_C1A0 16'hBBF1
`define CUBE_LUT_C1A1 16'hBBF1
`define CUBE_LUT_C1A2 16'hBBF1
`define CUBE_LUT_C1A3 16'hBBF1
`define CUBE_LUT_C1A4 16'hBBF2
`define CUBE_LUT_C1A5 16'hBBF2
`define CUBE_LUT_C1A6 16'hBBF2
`define CUBE_LUT_C1A7 16'hBBF2
`define CUBE_LUT_C1A8 16'hBBF2
`define CUBE_LUT_C1A9 16'hBBF2
`define CUBE_LUT_C1AA 16'hBBF2
`define CUBE_LUT_C1AB 16'hBBF2
`define CUBE_LUT_C1AC 16'hBBF2
`define CUBE_LUT_C1AD 16'hBBF2
`define CUBE_LUT_C1AE 16'hBBF2
`define CUBE_LUT_C1AF 16'hBBF2
`define CUBE_LUT_C1B0 16'hBBF2
`define CUBE_LUT_C1B1 16'hBBF2
`define CUBE_LUT_C1B2 16'hBBF2
`define CUBE_LUT_C1B3 16'hBBF2
`define CUBE_LUT_C1B4 16'hBBF2
`define CUBE_LUT_C1B5 16'hBBF2
`define CUBE_LUT_C1B6 16'hBBF2
`define CUBE_LUT_C1B7 16'hBBF3
`define CUBE_LUT_C1B8 16'hBBF3
`define CUBE_LUT_C1B9 16'hBBF3
`define CUBE_LUT_C1BA 16'hBBF3
`define CUBE_LUT_C1BB 16'hBBF3
`define CUBE_LUT_C1BC 16'hBBF3
`define CUBE_LUT_C1BD 16'hBBF3
`define CUBE_LUT_C1BE 16'hBBF3
`define CUBE_LUT_C1BF 16'hBBF3
`define CUBE_LUT_C1C0 16'hBBF3
`define CUBE_LUT_C1C1 16'hBBF3
`define CUBE_LUT_C1C2 16'hBBF3
`define CUBE_LUT_C1C3 16'hBBF3
`define CUBE_LUT_C1C4 16'hBBF3
`define CUBE_LUT_C1C5 16'hBBF3
`define CUBE_LUT_C1C6 16'hBBF3
`define CUBE_LUT_C1C7 16'hBBF3
`define CUBE_LUT_C1C8 16'hBBF3
`define CUBE_LUT_C1C9 16'hBBF3
`define CUBE_LUT_C1CA 16'hBBF4
`define CUBE_LUT_C1CB 16'hBBF4
`define CUBE_LUT_C1CC 16'hBBF4
`define CUBE_LUT_C1CD 16'hBBF4
`define CUBE_LUT_C1CE 16'hBBF4
`define CUBE_LUT_C1CF 16'hBBF4
`define CUBE_LUT_C1D0 16'hBBF4
`define CUBE_LUT_C1D1 16'hBBF4
`define CUBE_LUT_C1D2 16'hBBF4
`define CUBE_LUT_C1D3 16'hBBF4
`define CUBE_LUT_C1D4 16'hBBF4
`define CUBE_LUT_C1D5 16'hBBF4
`define CUBE_LUT_C1D6 16'hBBF4
`define CUBE_LUT_C1D7 16'hBBF4
`define CUBE_LUT_C1D8 16'hBBF4
`define CUBE_LUT_C1D9 16'hBBF4
`define CUBE_LUT_C1DA 16'hBBF4
`define CUBE_LUT_C1DB 16'hBBF4
`define CUBE_LUT_C1DC 16'hBBF4
`define CUBE_LUT_C1DD 16'hBBF4
`define CUBE_LUT_C1DE 16'hBBF4
`define CUBE_LUT_C1DF 16'hBBF4
`define CUBE_LUT_C1E0 16'hBBF5
`define CUBE_LUT_C1E1 16'hBBF5
`define CUBE_LUT_C1E2 16'hBBF5
`define CUBE_LUT_C1E3 16'hBBF5
`define CUBE_LUT_C1E4 16'hBBF5
`define CUBE_LUT_C1E5 16'hBBF5
`define CUBE_LUT_C1E6 16'hBBF5
`define CUBE_LUT_C1E7 16'hBBF5
`define CUBE_LUT_C1E8 16'hBBF5
`define CUBE_LUT_C1E9 16'hBBF5
`define CUBE_LUT_C1EA 16'hBBF5
`define CUBE_LUT_C1EB 16'hBBF5
`define CUBE_LUT_C1EC 16'hBBF5
`define CUBE_LUT_C1ED 16'hBBF5
`define CUBE_LUT_C1EE 16'hBBF5
`define CUBE_LUT_C1EF 16'hBBF5
`define CUBE_LUT_C1F0 16'hBBF5
`define CUBE_LUT_C1F1 16'hBBF5
`define CUBE_LUT_C1F2 16'hBBF5
`define CUBE_LUT_C1F3 16'hBBF5
`define CUBE_LUT_C1F4 16'hBBF5
`define CUBE_LUT_C1F5 16'hBBF5
`define CUBE_LUT_C1F6 16'hBBF5
`define CUBE_LUT_C1F7 16'hBBF6
`define CUBE_LUT_C1F8 16'hBBF6
`define CUBE_LUT_C1F9 16'hBBF6
`define CUBE_LUT_C1FA 16'hBBF6
`define CUBE_LUT_C1FB 16'hBBF6
`define CUBE_LUT_C1FC 16'hBBF6
`define CUBE_LUT_C1FD 16'hBBF6
`define CUBE_LUT_C1FE 16'hBBF6
`define CUBE_LUT_C1FF 16'hBBF6
`define CUBE_LUT_C200 16'hBBF6
