`define FP16_TO_INDEX_C200 0
`define FP16_TO_INDEX_C1FF 1
`define FP16_TO_INDEX_C1FE 2
`define FP16_TO_INDEX_C1FD 3
`define FP16_TO_INDEX_C1FC 4
`define FP16_TO_INDEX_C1FB 5
`define FP16_TO_INDEX_C1FA 6
`define FP16_TO_INDEX_C1F9 7
`define FP16_TO_INDEX_C1F8 8
`define FP16_TO_INDEX_C1F7 9
`define FP16_TO_INDEX_C1F6 10
`define FP16_TO_INDEX_C1F5 11
`define FP16_TO_INDEX_C1F4 12
`define FP16_TO_INDEX_C1F3 13
`define FP16_TO_INDEX_C1F2 14
`define FP16_TO_INDEX_C1F1 15
`define FP16_TO_INDEX_C1F0 16
`define FP16_TO_INDEX_C1EF 17
`define FP16_TO_INDEX_C1ED 18
`define FP16_TO_INDEX_C1EC 19
`define FP16_TO_INDEX_C1EB 20
`define FP16_TO_INDEX_C1EA 21
`define FP16_TO_INDEX_C1E9 22
`define FP16_TO_INDEX_C1E8 23
`define FP16_TO_INDEX_C1E7 24
`define FP16_TO_INDEX_C1E6 25
`define FP16_TO_INDEX_C1E5 26
`define FP16_TO_INDEX_C1E4 27
`define FP16_TO_INDEX_C1E3 28
`define FP16_TO_INDEX_C1E2 29
`define FP16_TO_INDEX_C1E1 30
`define FP16_TO_INDEX_C1E0 31
`define FP16_TO_INDEX_C1DF 32
`define FP16_TO_INDEX_C1DE 33
`define FP16_TO_INDEX_C1DD 34
`define FP16_TO_INDEX_C1DC 35
`define FP16_TO_INDEX_C1DB 36
`define FP16_TO_INDEX_C1DA 37
`define FP16_TO_INDEX_C1D9 38
`define FP16_TO_INDEX_C1D8 39
`define FP16_TO_INDEX_C1D7 40
`define FP16_TO_INDEX_C1D6 41
`define FP16_TO_INDEX_C1D5 42
`define FP16_TO_INDEX_C1D4 43
`define FP16_TO_INDEX_C1D3 44
`define FP16_TO_INDEX_C1D2 45
`define FP16_TO_INDEX_C1D1 46
`define FP16_TO_INDEX_C1D0 47
`define FP16_TO_INDEX_C1CF 48
`define FP16_TO_INDEX_C1CE 49
`define FP16_TO_INDEX_C1CD 50
`define FP16_TO_INDEX_C1CC 51
`define FP16_TO_INDEX_C1CB 52
`define FP16_TO_INDEX_C1C9 53
`define FP16_TO_INDEX_C1C8 54
`define FP16_TO_INDEX_C1C7 55
`define FP16_TO_INDEX_C1C6 56
`define FP16_TO_INDEX_C1C5 57
`define FP16_TO_INDEX_C1C4 58
`define FP16_TO_INDEX_C1C3 59
`define FP16_TO_INDEX_C1C2 60
`define FP16_TO_INDEX_C1C1 61
`define FP16_TO_INDEX_C1C0 62
`define FP16_TO_INDEX_C1BF 63
`define FP16_TO_INDEX_C1BE 64
`define FP16_TO_INDEX_C1BD 65
`define FP16_TO_INDEX_C1BC 66
`define FP16_TO_INDEX_C1BB 67
`define FP16_TO_INDEX_C1BA 68
`define FP16_TO_INDEX_C1B9 69
`define FP16_TO_INDEX_C1B8 70
`define FP16_TO_INDEX_C1B7 71
`define FP16_TO_INDEX_C1B6 72
`define FP16_TO_INDEX_C1B5 73
`define FP16_TO_INDEX_C1B4 74
`define FP16_TO_INDEX_C1B3 75
`define FP16_TO_INDEX_C1B2 76
`define FP16_TO_INDEX_C1B1 77
`define FP16_TO_INDEX_C1B0 78
`define FP16_TO_INDEX_C1AF 79
`define FP16_TO_INDEX_C1AE 80
`define FP16_TO_INDEX_C1AD 81
`define FP16_TO_INDEX_C1AC 82
`define FP16_TO_INDEX_C1AB 83
`define FP16_TO_INDEX_C1AA 84
`define FP16_TO_INDEX_C1A9 85
`define FP16_TO_INDEX_C1A8 86
`define FP16_TO_INDEX_C1A7 87
`define FP16_TO_INDEX_C1A5 88
`define FP16_TO_INDEX_C1A4 89
`define FP16_TO_INDEX_C1A3 90
`define FP16_TO_INDEX_C1A2 91
`define FP16_TO_INDEX_C1A1 92
`define FP16_TO_INDEX_C1A0 93
`define FP16_TO_INDEX_C19F 94
`define FP16_TO_INDEX_C19E 95
`define FP16_TO_INDEX_C19D 96
`define FP16_TO_INDEX_C19C 97
`define FP16_TO_INDEX_C19B 98
`define FP16_TO_INDEX_C19A 99
`define FP16_TO_INDEX_C199 100
`define FP16_TO_INDEX_C198 101
`define FP16_TO_INDEX_C197 102
`define FP16_TO_INDEX_C196 103
`define FP16_TO_INDEX_C195 104
`define FP16_TO_INDEX_C194 105
`define FP16_TO_INDEX_C193 106
`define FP16_TO_INDEX_C192 107
`define FP16_TO_INDEX_C191 108
`define FP16_TO_INDEX_C190 109
`define FP16_TO_INDEX_C18F 110
`define FP16_TO_INDEX_C18E 111
`define FP16_TO_INDEX_C18D 112
`define FP16_TO_INDEX_C18C 113
`define FP16_TO_INDEX_C18B 114
`define FP16_TO_INDEX_C18A 115
`define FP16_TO_INDEX_C189 116
`define FP16_TO_INDEX_C188 117
`define FP16_TO_INDEX_C187 118
`define FP16_TO_INDEX_C186 119
`define FP16_TO_INDEX_C185 120
`define FP16_TO_INDEX_C184 121
`define FP16_TO_INDEX_C183 122
`define FP16_TO_INDEX_C181 123
`define FP16_TO_INDEX_C180 124
`define FP16_TO_INDEX_C17F 125
`define FP16_TO_INDEX_C17E 126
`define FP16_TO_INDEX_C17D 127
`define FP16_TO_INDEX_C17C 128
`define FP16_TO_INDEX_C17B 129
`define FP16_TO_INDEX_C17A 130
`define FP16_TO_INDEX_C179 131
`define FP16_TO_INDEX_C178 132
`define FP16_TO_INDEX_C177 133
`define FP16_TO_INDEX_C176 134
`define FP16_TO_INDEX_C175 135
`define FP16_TO_INDEX_C174 136
`define FP16_TO_INDEX_C173 137
`define FP16_TO_INDEX_C172 138
`define FP16_TO_INDEX_C171 139
`define FP16_TO_INDEX_C170 140
`define FP16_TO_INDEX_C16F 141
`define FP16_TO_INDEX_C16E 142
`define FP16_TO_INDEX_C16D 143
`define FP16_TO_INDEX_C16C 144
`define FP16_TO_INDEX_C16B 145
`define FP16_TO_INDEX_C16A 146
`define FP16_TO_INDEX_C169 147
`define FP16_TO_INDEX_C168 148
`define FP16_TO_INDEX_C167 149
`define FP16_TO_INDEX_C166 150
`define FP16_TO_INDEX_C165 151
`define FP16_TO_INDEX_C164 152
`define FP16_TO_INDEX_C163 153
`define FP16_TO_INDEX_C162 154
`define FP16_TO_INDEX_C161 155
`define FP16_TO_INDEX_C160 156
`define FP16_TO_INDEX_C15F 157
`define FP16_TO_INDEX_C15E 158
`define FP16_TO_INDEX_C15C 159
`define FP16_TO_INDEX_C15B 160
`define FP16_TO_INDEX_C15A 161
`define FP16_TO_INDEX_C159 162
`define FP16_TO_INDEX_C158 163
`define FP16_TO_INDEX_C157 164
`define FP16_TO_INDEX_C156 165
`define FP16_TO_INDEX_C155 166
`define FP16_TO_INDEX_C154 167
`define FP16_TO_INDEX_C153 168
`define FP16_TO_INDEX_C152 169
`define FP16_TO_INDEX_C151 170
`define FP16_TO_INDEX_C150 171
`define FP16_TO_INDEX_C14F 172
`define FP16_TO_INDEX_C14E 173
`define FP16_TO_INDEX_C14D 174
`define FP16_TO_INDEX_C14C 175
`define FP16_TO_INDEX_C14B 176
`define FP16_TO_INDEX_C14A 177
`define FP16_TO_INDEX_C149 178
`define FP16_TO_INDEX_C148 179
`define FP16_TO_INDEX_C147 180
`define FP16_TO_INDEX_C146 181
`define FP16_TO_INDEX_C145 182
`define FP16_TO_INDEX_C144 183
`define FP16_TO_INDEX_C143 184
`define FP16_TO_INDEX_C142 185
`define FP16_TO_INDEX_C141 186
`define FP16_TO_INDEX_C140 187
`define FP16_TO_INDEX_C13F 188
`define FP16_TO_INDEX_C13E 189
`define FP16_TO_INDEX_C13D 190
`define FP16_TO_INDEX_C13C 191
`define FP16_TO_INDEX_C13B 192
`define FP16_TO_INDEX_C13A 193
`define FP16_TO_INDEX_C138 194
`define FP16_TO_INDEX_C137 195
`define FP16_TO_INDEX_C136 196
`define FP16_TO_INDEX_C135 197
`define FP16_TO_INDEX_C134 198
`define FP16_TO_INDEX_C133 199
`define FP16_TO_INDEX_C132 200
`define FP16_TO_INDEX_C131 201
`define FP16_TO_INDEX_C130 202
`define FP16_TO_INDEX_C12F 203
`define FP16_TO_INDEX_C12E 204
`define FP16_TO_INDEX_C12D 205
`define FP16_TO_INDEX_C12C 206
`define FP16_TO_INDEX_C12B 207
`define FP16_TO_INDEX_C12A 208
`define FP16_TO_INDEX_C129 209
`define FP16_TO_INDEX_C128 210
`define FP16_TO_INDEX_C127 211
`define FP16_TO_INDEX_C126 212
`define FP16_TO_INDEX_C125 213
`define FP16_TO_INDEX_C124 214
`define FP16_TO_INDEX_C123 215
`define FP16_TO_INDEX_C122 216
`define FP16_TO_INDEX_C121 217
`define FP16_TO_INDEX_C120 218
`define FP16_TO_INDEX_C11F 219
`define FP16_TO_INDEX_C11E 220
`define FP16_TO_INDEX_C11D 221
`define FP16_TO_INDEX_C11C 222
`define FP16_TO_INDEX_C11B 223
`define FP16_TO_INDEX_C11A 224
`define FP16_TO_INDEX_C119 225
`define FP16_TO_INDEX_C118 226
`define FP16_TO_INDEX_C117 227
`define FP16_TO_INDEX_C116 228
`define FP16_TO_INDEX_C114 229
`define FP16_TO_INDEX_C113 230
`define FP16_TO_INDEX_C112 231
`define FP16_TO_INDEX_C111 232
`define FP16_TO_INDEX_C110 233
`define FP16_TO_INDEX_C10F 234
`define FP16_TO_INDEX_C10E 235
`define FP16_TO_INDEX_C10D 236
`define FP16_TO_INDEX_C10C 237
`define FP16_TO_INDEX_C10B 238
`define FP16_TO_INDEX_C10A 239
`define FP16_TO_INDEX_C109 240
`define FP16_TO_INDEX_C108 241
`define FP16_TO_INDEX_C107 242
`define FP16_TO_INDEX_C106 243
`define FP16_TO_INDEX_C105 244
`define FP16_TO_INDEX_C104 245
`define FP16_TO_INDEX_C103 246
`define FP16_TO_INDEX_C102 247
`define FP16_TO_INDEX_C101 248
`define FP16_TO_INDEX_C100 249
`define FP16_TO_INDEX_C0FF 250
`define FP16_TO_INDEX_C0FE 251
`define FP16_TO_INDEX_C0FD 252
`define FP16_TO_INDEX_C0FC 253
`define FP16_TO_INDEX_C0FB 254
`define FP16_TO_INDEX_C0FA 255
`define FP16_TO_INDEX_C0F9 256
`define FP16_TO_INDEX_C0F8 257
`define FP16_TO_INDEX_C0F7 258
`define FP16_TO_INDEX_C0F6 259
`define FP16_TO_INDEX_C0F5 260
`define FP16_TO_INDEX_C0F4 261
`define FP16_TO_INDEX_C0F3 262
`define FP16_TO_INDEX_C0F2 263
`define FP16_TO_INDEX_C0F0 264
`define FP16_TO_INDEX_C0EF 265
`define FP16_TO_INDEX_C0EE 266
`define FP16_TO_INDEX_C0ED 267
`define FP16_TO_INDEX_C0EC 268
`define FP16_TO_INDEX_C0EB 269
`define FP16_TO_INDEX_C0EA 270
`define FP16_TO_INDEX_C0E9 271
`define FP16_TO_INDEX_C0E8 272
`define FP16_TO_INDEX_C0E7 273
`define FP16_TO_INDEX_C0E6 274
`define FP16_TO_INDEX_C0E5 275
`define FP16_TO_INDEX_C0E4 276
`define FP16_TO_INDEX_C0E3 277
`define FP16_TO_INDEX_C0E2 278
`define FP16_TO_INDEX_C0E1 279
`define FP16_TO_INDEX_C0E0 280
`define FP16_TO_INDEX_C0DF 281
`define FP16_TO_INDEX_C0DE 282
`define FP16_TO_INDEX_C0DD 283
`define FP16_TO_INDEX_C0DC 284
`define FP16_TO_INDEX_C0DB 285
`define FP16_TO_INDEX_C0DA 286
`define FP16_TO_INDEX_C0D9 287
`define FP16_TO_INDEX_C0D8 288
`define FP16_TO_INDEX_C0D7 289
`define FP16_TO_INDEX_C0D6 290
`define FP16_TO_INDEX_C0D5 291
`define FP16_TO_INDEX_C0D4 292
`define FP16_TO_INDEX_C0D3 293
`define FP16_TO_INDEX_C0D2 294
`define FP16_TO_INDEX_C0D1 295
`define FP16_TO_INDEX_C0D0 296
`define FP16_TO_INDEX_C0CF 297
`define FP16_TO_INDEX_C0CE 298
`define FP16_TO_INDEX_C0CC 299
`define FP16_TO_INDEX_C0CB 300
`define FP16_TO_INDEX_C0CA 301
`define FP16_TO_INDEX_C0C9 302
`define FP16_TO_INDEX_C0C8 303
`define FP16_TO_INDEX_C0C7 304
`define FP16_TO_INDEX_C0C6 305
`define FP16_TO_INDEX_C0C5 306
`define FP16_TO_INDEX_C0C4 307
`define FP16_TO_INDEX_C0C3 308
`define FP16_TO_INDEX_C0C2 309
`define FP16_TO_INDEX_C0C1 310
`define FP16_TO_INDEX_C0C0 311
`define FP16_TO_INDEX_C0BF 312
`define FP16_TO_INDEX_C0BE 313
`define FP16_TO_INDEX_C0BD 314
`define FP16_TO_INDEX_C0BC 315
`define FP16_TO_INDEX_C0BB 316
`define FP16_TO_INDEX_C0BA 317
`define FP16_TO_INDEX_C0B9 318
`define FP16_TO_INDEX_C0B8 319
`define FP16_TO_INDEX_C0B7 320
`define FP16_TO_INDEX_C0B6 321
`define FP16_TO_INDEX_C0B5 322
`define FP16_TO_INDEX_C0B4 323
`define FP16_TO_INDEX_C0B3 324
`define FP16_TO_INDEX_C0B2 325
`define FP16_TO_INDEX_C0B1 326
`define FP16_TO_INDEX_C0B0 327
`define FP16_TO_INDEX_C0AF 328
`define FP16_TO_INDEX_C0AE 329
`define FP16_TO_INDEX_C0AD 330
`define FP16_TO_INDEX_C0AC 331
`define FP16_TO_INDEX_C0AB 332
`define FP16_TO_INDEX_C0AA 333
`define FP16_TO_INDEX_C0A8 334
`define FP16_TO_INDEX_C0A7 335
`define FP16_TO_INDEX_C0A6 336
`define FP16_TO_INDEX_C0A5 337
`define FP16_TO_INDEX_C0A4 338
`define FP16_TO_INDEX_C0A3 339
`define FP16_TO_INDEX_C0A2 340
`define FP16_TO_INDEX_C0A1 341
`define FP16_TO_INDEX_C0A0 342
`define FP16_TO_INDEX_C09F 343
`define FP16_TO_INDEX_C09E 344
`define FP16_TO_INDEX_C09D 345
`define FP16_TO_INDEX_C09C 346
`define FP16_TO_INDEX_C09B 347
`define FP16_TO_INDEX_C09A 348
`define FP16_TO_INDEX_C099 349
`define FP16_TO_INDEX_C098 350
`define FP16_TO_INDEX_C097 351
`define FP16_TO_INDEX_C096 352
`define FP16_TO_INDEX_C095 353
`define FP16_TO_INDEX_C094 354
`define FP16_TO_INDEX_C093 355
`define FP16_TO_INDEX_C092 356
`define FP16_TO_INDEX_C091 357
`define FP16_TO_INDEX_C090 358
`define FP16_TO_INDEX_C08F 359
`define FP16_TO_INDEX_C08E 360
`define FP16_TO_INDEX_C08D 361
`define FP16_TO_INDEX_C08C 362
`define FP16_TO_INDEX_C08B 363
`define FP16_TO_INDEX_C08A 364
`define FP16_TO_INDEX_C089 365
`define FP16_TO_INDEX_C088 366
`define FP16_TO_INDEX_C087 367
`define FP16_TO_INDEX_C086 368
`define FP16_TO_INDEX_C084 369
`define FP16_TO_INDEX_C083 370
`define FP16_TO_INDEX_C082 371
`define FP16_TO_INDEX_C081 372
`define FP16_TO_INDEX_C080 373
`define FP16_TO_INDEX_C07F 374
`define FP16_TO_INDEX_C07E 375
`define FP16_TO_INDEX_C07D 376
`define FP16_TO_INDEX_C07C 377
`define FP16_TO_INDEX_C07B 378
`define FP16_TO_INDEX_C07A 379
`define FP16_TO_INDEX_C079 380
`define FP16_TO_INDEX_C078 381
`define FP16_TO_INDEX_C077 382
`define FP16_TO_INDEX_C076 383
`define FP16_TO_INDEX_C075 384
`define FP16_TO_INDEX_C074 385
`define FP16_TO_INDEX_C073 386
`define FP16_TO_INDEX_C072 387
`define FP16_TO_INDEX_C071 388
`define FP16_TO_INDEX_C070 389
`define FP16_TO_INDEX_C06F 390
`define FP16_TO_INDEX_C06E 391
`define FP16_TO_INDEX_C06D 392
`define FP16_TO_INDEX_C06C 393
`define FP16_TO_INDEX_C06B 394
`define FP16_TO_INDEX_C06A 395
`define FP16_TO_INDEX_C069 396
`define FP16_TO_INDEX_C068 397
`define FP16_TO_INDEX_C067 398
`define FP16_TO_INDEX_C066 399
`define FP16_TO_INDEX_C065 400
`define FP16_TO_INDEX_C064 401
`define FP16_TO_INDEX_C063 402
`define FP16_TO_INDEX_C062 403
`define FP16_TO_INDEX_C061 404
`define FP16_TO_INDEX_C05F 405
`define FP16_TO_INDEX_C05E 406
`define FP16_TO_INDEX_C05D 407
`define FP16_TO_INDEX_C05C 408
`define FP16_TO_INDEX_C05B 409
`define FP16_TO_INDEX_C05A 410
`define FP16_TO_INDEX_C059 411
`define FP16_TO_INDEX_C058 412
`define FP16_TO_INDEX_C057 413
`define FP16_TO_INDEX_C056 414
`define FP16_TO_INDEX_C055 415
`define FP16_TO_INDEX_C054 416
`define FP16_TO_INDEX_C053 417
`define FP16_TO_INDEX_C052 418
`define FP16_TO_INDEX_C051 419
`define FP16_TO_INDEX_C050 420
`define FP16_TO_INDEX_C04F 421
`define FP16_TO_INDEX_C04E 422
`define FP16_TO_INDEX_C04D 423
`define FP16_TO_INDEX_C04C 424
`define FP16_TO_INDEX_C04B 425
`define FP16_TO_INDEX_C04A 426
`define FP16_TO_INDEX_C049 427
`define FP16_TO_INDEX_C048 428
`define FP16_TO_INDEX_C047 429
`define FP16_TO_INDEX_C046 430
`define FP16_TO_INDEX_C045 431
`define FP16_TO_INDEX_C044 432
`define FP16_TO_INDEX_C043 433
`define FP16_TO_INDEX_C042 434
`define FP16_TO_INDEX_C041 435
`define FP16_TO_INDEX_C040 436
`define FP16_TO_INDEX_C03F 437
`define FP16_TO_INDEX_C03E 438
`define FP16_TO_INDEX_C03D 439
`define FP16_TO_INDEX_C03B 440
`define FP16_TO_INDEX_C03A 441
`define FP16_TO_INDEX_C039 442
`define FP16_TO_INDEX_C038 443
`define FP16_TO_INDEX_C037 444
`define FP16_TO_INDEX_C036 445
`define FP16_TO_INDEX_C035 446
`define FP16_TO_INDEX_C034 447
`define FP16_TO_INDEX_C033 448
`define FP16_TO_INDEX_C032 449
`define FP16_TO_INDEX_C031 450
`define FP16_TO_INDEX_C030 451
`define FP16_TO_INDEX_C02F 452
`define FP16_TO_INDEX_C02E 453
`define FP16_TO_INDEX_C02D 454
`define FP16_TO_INDEX_C02C 455
`define FP16_TO_INDEX_C02B 456
`define FP16_TO_INDEX_C02A 457
`define FP16_TO_INDEX_C029 458
`define FP16_TO_INDEX_C028 459
`define FP16_TO_INDEX_C027 460
`define FP16_TO_INDEX_C026 461
`define FP16_TO_INDEX_C025 462
`define FP16_TO_INDEX_C024 463
`define FP16_TO_INDEX_C023 464
`define FP16_TO_INDEX_C022 465
`define FP16_TO_INDEX_C021 466
`define FP16_TO_INDEX_C020 467
`define FP16_TO_INDEX_C01F 468
`define FP16_TO_INDEX_C01E 469
`define FP16_TO_INDEX_C01D 470
`define FP16_TO_INDEX_C01C 471
`define FP16_TO_INDEX_C01B 472
`define FP16_TO_INDEX_C01A 473
`define FP16_TO_INDEX_C019 474
`define FP16_TO_INDEX_C017 475
`define FP16_TO_INDEX_C016 476
`define FP16_TO_INDEX_C015 477
`define FP16_TO_INDEX_C014 478
`define FP16_TO_INDEX_C013 479
`define FP16_TO_INDEX_C012 480
`define FP16_TO_INDEX_C011 481
`define FP16_TO_INDEX_C010 482
`define FP16_TO_INDEX_C00F 483
`define FP16_TO_INDEX_C00E 484
`define FP16_TO_INDEX_C00D 485
`define FP16_TO_INDEX_C00C 486
`define FP16_TO_INDEX_C00B 487
`define FP16_TO_INDEX_C00A 488
`define FP16_TO_INDEX_C009 489
`define FP16_TO_INDEX_C008 490
`define FP16_TO_INDEX_C007 491
`define FP16_TO_INDEX_C006 492
`define FP16_TO_INDEX_C005 493
`define FP16_TO_INDEX_C004 494
`define FP16_TO_INDEX_C003 495
`define FP16_TO_INDEX_C002 496
`define FP16_TO_INDEX_C001 497
`define FP16_TO_INDEX_C000 498
`define FP16_TO_INDEX_BFFE 499
`define FP16_TO_INDEX_BFFC 500
`define FP16_TO_INDEX_BFF9 501
`define FP16_TO_INDEX_BFF7 502
`define FP16_TO_INDEX_BFF5 503
`define FP16_TO_INDEX_BFF3 504
`define FP16_TO_INDEX_BFF1 505
`define FP16_TO_INDEX_BFEF 506
`define FP16_TO_INDEX_BFED 507
`define FP16_TO_INDEX_BFEB 508
`define FP16_TO_INDEX_BFE9 509
`define FP16_TO_INDEX_BFE7 510
`define FP16_TO_INDEX_BFE5 511
`define FP16_TO_INDEX_BFE3 512
`define FP16_TO_INDEX_BFE1 513
`define FP16_TO_INDEX_BFDF 514
`define FP16_TO_INDEX_BFDD 515
`define FP16_TO_INDEX_BFDB 516
`define FP16_TO_INDEX_BFD9 517
`define FP16_TO_INDEX_BFD7 518
`define FP16_TO_INDEX_BFD4 519
`define FP16_TO_INDEX_BFD2 520
`define FP16_TO_INDEX_BFD0 521
`define FP16_TO_INDEX_BFCE 522
`define FP16_TO_INDEX_BFCC 523
`define FP16_TO_INDEX_BFCA 524
`define FP16_TO_INDEX_BFC8 525
`define FP16_TO_INDEX_BFC6 526
`define FP16_TO_INDEX_BFC4 527
`define FP16_TO_INDEX_BFC2 528
`define FP16_TO_INDEX_BFC0 529
`define FP16_TO_INDEX_BFBE 530
`define FP16_TO_INDEX_BFBC 531
`define FP16_TO_INDEX_BFBA 532
`define FP16_TO_INDEX_BFB8 533
`define FP16_TO_INDEX_BFB6 534
`define FP16_TO_INDEX_BFB4 535
`define FP16_TO_INDEX_BFB1 536
`define FP16_TO_INDEX_BFAF 537
`define FP16_TO_INDEX_BFAD 538
`define FP16_TO_INDEX_BFAB 539
`define FP16_TO_INDEX_BFA9 540
`define FP16_TO_INDEX_BFA7 541
`define FP16_TO_INDEX_BFA5 542
`define FP16_TO_INDEX_BFA3 543
`define FP16_TO_INDEX_BFA1 544
`define FP16_TO_INDEX_BF9F 545
`define FP16_TO_INDEX_BF9D 546
`define FP16_TO_INDEX_BF9B 547
`define FP16_TO_INDEX_BF99 548
`define FP16_TO_INDEX_BF97 549
`define FP16_TO_INDEX_BF95 550
`define FP16_TO_INDEX_BF93 551
`define FP16_TO_INDEX_BF91 552
`define FP16_TO_INDEX_BF8F 553
`define FP16_TO_INDEX_BF8C 554
`define FP16_TO_INDEX_BF8A 555
`define FP16_TO_INDEX_BF88 556
`define FP16_TO_INDEX_BF86 557
`define FP16_TO_INDEX_BF84 558
`define FP16_TO_INDEX_BF82 559
`define FP16_TO_INDEX_BF80 560
`define FP16_TO_INDEX_BF7E 561
`define FP16_TO_INDEX_BF7C 562
`define FP16_TO_INDEX_BF7A 563
`define FP16_TO_INDEX_BF78 564
`define FP16_TO_INDEX_BF76 565
`define FP16_TO_INDEX_BF74 566
`define FP16_TO_INDEX_BF72 567
`define FP16_TO_INDEX_BF70 568
`define FP16_TO_INDEX_BF6E 569
`define FP16_TO_INDEX_BF6C 570
`define FP16_TO_INDEX_BF6A 571
`define FP16_TO_INDEX_BF67 572
`define FP16_TO_INDEX_BF65 573
`define FP16_TO_INDEX_BF63 574
`define FP16_TO_INDEX_BF61 575
`define FP16_TO_INDEX_BF5F 576
`define FP16_TO_INDEX_BF5D 577
`define FP16_TO_INDEX_BF5B 578
`define FP16_TO_INDEX_BF59 579
`define FP16_TO_INDEX_BF57 580
`define FP16_TO_INDEX_BF55 581
`define FP16_TO_INDEX_BF53 582
`define FP16_TO_INDEX_BF51 583
`define FP16_TO_INDEX_BF4F 584
`define FP16_TO_INDEX_BF4D 585
`define FP16_TO_INDEX_BF4B 586
`define FP16_TO_INDEX_BF49 587
`define FP16_TO_INDEX_BF47 588
`define FP16_TO_INDEX_BF44 589
`define FP16_TO_INDEX_BF42 590
`define FP16_TO_INDEX_BF40 591
`define FP16_TO_INDEX_BF3E 592
`define FP16_TO_INDEX_BF3C 593
`define FP16_TO_INDEX_BF3A 594
`define FP16_TO_INDEX_BF38 595
`define FP16_TO_INDEX_BF36 596
`define FP16_TO_INDEX_BF34 597
`define FP16_TO_INDEX_BF32 598
`define FP16_TO_INDEX_BF30 599
`define FP16_TO_INDEX_BF2E 600
`define FP16_TO_INDEX_BF2C 601
`define FP16_TO_INDEX_BF2A 602
`define FP16_TO_INDEX_BF28 603
`define FP16_TO_INDEX_BF26 604
`define FP16_TO_INDEX_BF24 605
`define FP16_TO_INDEX_BF22 606
`define FP16_TO_INDEX_BF1F 607
`define FP16_TO_INDEX_BF1D 608
`define FP16_TO_INDEX_BF1B 609
`define FP16_TO_INDEX_BF19 610
`define FP16_TO_INDEX_BF17 611
`define FP16_TO_INDEX_BF15 612
`define FP16_TO_INDEX_BF13 613
`define FP16_TO_INDEX_BF11 614
`define FP16_TO_INDEX_BF0F 615
`define FP16_TO_INDEX_BF0D 616
`define FP16_TO_INDEX_BF0B 617
`define FP16_TO_INDEX_BF09 618
`define FP16_TO_INDEX_BF07 619
`define FP16_TO_INDEX_BF05 620
`define FP16_TO_INDEX_BF03 621
`define FP16_TO_INDEX_BF01 622
`define FP16_TO_INDEX_BEFF 623
`define FP16_TO_INDEX_BEFC 624
`define FP16_TO_INDEX_BEFA 625
`define FP16_TO_INDEX_BEF8 626
`define FP16_TO_INDEX_BEF6 627
`define FP16_TO_INDEX_BEF4 628
`define FP16_TO_INDEX_BEF2 629
`define FP16_TO_INDEX_BEF0 630
`define FP16_TO_INDEX_BEEE 631
`define FP16_TO_INDEX_BEEC 632
`define FP16_TO_INDEX_BEEA 633
`define FP16_TO_INDEX_BEE8 634
`define FP16_TO_INDEX_BEE6 635
`define FP16_TO_INDEX_BEE4 636
`define FP16_TO_INDEX_BEE2 637
`define FP16_TO_INDEX_BEE0 638
`define FP16_TO_INDEX_BEDE 639
`define FP16_TO_INDEX_BEDC 640
`define FP16_TO_INDEX_BEDA 641
`define FP16_TO_INDEX_BED7 642
`define FP16_TO_INDEX_BED5 643
`define FP16_TO_INDEX_BED3 644
`define FP16_TO_INDEX_BED1 645
`define FP16_TO_INDEX_BECF 646
`define FP16_TO_INDEX_BECD 647
`define FP16_TO_INDEX_BECB 648
`define FP16_TO_INDEX_BEC9 649
`define FP16_TO_INDEX_BEC7 650
`define FP16_TO_INDEX_BEC5 651
`define FP16_TO_INDEX_BEC3 652
`define FP16_TO_INDEX_BEC1 653
`define FP16_TO_INDEX_BEBF 654
`define FP16_TO_INDEX_BEBD 655
`define FP16_TO_INDEX_BEBB 656
`define FP16_TO_INDEX_BEB9 657
`define FP16_TO_INDEX_BEB7 658
`define FP16_TO_INDEX_BEB4 659
`define FP16_TO_INDEX_BEB2 660
`define FP16_TO_INDEX_BEB0 661
`define FP16_TO_INDEX_BEAE 662
`define FP16_TO_INDEX_BEAC 663
`define FP16_TO_INDEX_BEAA 664
`define FP16_TO_INDEX_BEA8 665
`define FP16_TO_INDEX_BEA6 666
`define FP16_TO_INDEX_BEA4 667
`define FP16_TO_INDEX_BEA2 668
`define FP16_TO_INDEX_BEA0 669
`define FP16_TO_INDEX_BE9E 670
`define FP16_TO_INDEX_BE9C 671
`define FP16_TO_INDEX_BE9A 672
`define FP16_TO_INDEX_BE98 673
`define FP16_TO_INDEX_BE96 674
`define FP16_TO_INDEX_BE94 675
`define FP16_TO_INDEX_BE92 676
`define FP16_TO_INDEX_BE8F 677
`define FP16_TO_INDEX_BE8D 678
`define FP16_TO_INDEX_BE8B 679
`define FP16_TO_INDEX_BE89 680
`define FP16_TO_INDEX_BE87 681
`define FP16_TO_INDEX_BE85 682
`define FP16_TO_INDEX_BE83 683
`define FP16_TO_INDEX_BE81 684
`define FP16_TO_INDEX_BE7F 685
`define FP16_TO_INDEX_BE7D 686
`define FP16_TO_INDEX_BE7B 687
`define FP16_TO_INDEX_BE79 688
`define FP16_TO_INDEX_BE77 689
`define FP16_TO_INDEX_BE75 690
`define FP16_TO_INDEX_BE73 691
`define FP16_TO_INDEX_BE71 692
`define FP16_TO_INDEX_BE6F 693
`define FP16_TO_INDEX_BE6D 694
`define FP16_TO_INDEX_BE6A 695
`define FP16_TO_INDEX_BE68 696
`define FP16_TO_INDEX_BE66 697
`define FP16_TO_INDEX_BE64 698
`define FP16_TO_INDEX_BE62 699
`define FP16_TO_INDEX_BE60 700
`define FP16_TO_INDEX_BE5E 701
`define FP16_TO_INDEX_BE5C 702
`define FP16_TO_INDEX_BE5A 703
`define FP16_TO_INDEX_BE58 704
`define FP16_TO_INDEX_BE56 705
`define FP16_TO_INDEX_BE54 706
`define FP16_TO_INDEX_BE52 707
`define FP16_TO_INDEX_BE50 708
`define FP16_TO_INDEX_BE4E 709
`define FP16_TO_INDEX_BE4C 710
`define FP16_TO_INDEX_BE4A 711
`define FP16_TO_INDEX_BE47 712
`define FP16_TO_INDEX_BE45 713
`define FP16_TO_INDEX_BE43 714
`define FP16_TO_INDEX_BE41 715
`define FP16_TO_INDEX_BE3F 716
`define FP16_TO_INDEX_BE3D 717
`define FP16_TO_INDEX_BE3B 718
`define FP16_TO_INDEX_BE39 719
`define FP16_TO_INDEX_BE37 720
`define FP16_TO_INDEX_BE35 721
`define FP16_TO_INDEX_BE33 722
`define FP16_TO_INDEX_BE31 723
`define FP16_TO_INDEX_BE2F 724
`define FP16_TO_INDEX_BE2D 725
`define FP16_TO_INDEX_BE2B 726
`define FP16_TO_INDEX_BE29 727
`define FP16_TO_INDEX_BE27 728
`define FP16_TO_INDEX_BE25 729
`define FP16_TO_INDEX_BE22 730
`define FP16_TO_INDEX_BE20 731
`define FP16_TO_INDEX_BE1E 732
`define FP16_TO_INDEX_BE1C 733
`define FP16_TO_INDEX_BE1A 734
`define FP16_TO_INDEX_BE18 735
`define FP16_TO_INDEX_BE16 736
`define FP16_TO_INDEX_BE14 737
`define FP16_TO_INDEX_BE12 738
`define FP16_TO_INDEX_BE10 739
`define FP16_TO_INDEX_BE0E 740
`define FP16_TO_INDEX_BE0C 741
`define FP16_TO_INDEX_BE0A 742
`define FP16_TO_INDEX_BE08 743
`define FP16_TO_INDEX_BE06 744
`define FP16_TO_INDEX_BE04 745
`define FP16_TO_INDEX_BE02 746
`define FP16_TO_INDEX_BDFF 747
`define FP16_TO_INDEX_BDFD 748
`define FP16_TO_INDEX_BDFB 749
`define FP16_TO_INDEX_BDF9 750
`define FP16_TO_INDEX_BDF7 751
`define FP16_TO_INDEX_BDF5 752
`define FP16_TO_INDEX_BDF3 753
`define FP16_TO_INDEX_BDF1 754
`define FP16_TO_INDEX_BDEF 755
`define FP16_TO_INDEX_BDED 756
`define FP16_TO_INDEX_BDEB 757
`define FP16_TO_INDEX_BDE9 758
`define FP16_TO_INDEX_BDE7 759
`define FP16_TO_INDEX_BDE5 760
`define FP16_TO_INDEX_BDE3 761
`define FP16_TO_INDEX_BDE1 762
`define FP16_TO_INDEX_BDDF 763
`define FP16_TO_INDEX_BDDD 764
`define FP16_TO_INDEX_BDDA 765
`define FP16_TO_INDEX_BDD8 766
`define FP16_TO_INDEX_BDD6 767
`define FP16_TO_INDEX_BDD4 768
`define FP16_TO_INDEX_BDD2 769
`define FP16_TO_INDEX_BDD0 770
`define FP16_TO_INDEX_BDCE 771
`define FP16_TO_INDEX_BDCC 772
`define FP16_TO_INDEX_BDCA 773
`define FP16_TO_INDEX_BDC8 774
`define FP16_TO_INDEX_BDC6 775
`define FP16_TO_INDEX_BDC4 776
`define FP16_TO_INDEX_BDC2 777
`define FP16_TO_INDEX_BDC0 778
`define FP16_TO_INDEX_BDBE 779
`define FP16_TO_INDEX_BDBC 780
`define FP16_TO_INDEX_BDBA 781
`define FP16_TO_INDEX_BDB7 782
`define FP16_TO_INDEX_BDB5 783
`define FP16_TO_INDEX_BDB3 784
`define FP16_TO_INDEX_BDB1 785
`define FP16_TO_INDEX_BDAF 786
`define FP16_TO_INDEX_BDAD 787
`define FP16_TO_INDEX_BDAB 788
`define FP16_TO_INDEX_BDA9 789
`define FP16_TO_INDEX_BDA7 790
`define FP16_TO_INDEX_BDA5 791
`define FP16_TO_INDEX_BDA3 792
`define FP16_TO_INDEX_BDA1 793
`define FP16_TO_INDEX_BD9F 794
`define FP16_TO_INDEX_BD9D 795
`define FP16_TO_INDEX_BD9B 796
`define FP16_TO_INDEX_BD99 797
`define FP16_TO_INDEX_BD97 798
`define FP16_TO_INDEX_BD95 799
`define FP16_TO_INDEX_BD92 800
`define FP16_TO_INDEX_BD90 801
`define FP16_TO_INDEX_BD8E 802
`define FP16_TO_INDEX_BD8C 803
`define FP16_TO_INDEX_BD8A 804
`define FP16_TO_INDEX_BD88 805
`define FP16_TO_INDEX_BD86 806
`define FP16_TO_INDEX_BD84 807
`define FP16_TO_INDEX_BD82 808
`define FP16_TO_INDEX_BD80 809
`define FP16_TO_INDEX_BD7E 810
`define FP16_TO_INDEX_BD7C 811
`define FP16_TO_INDEX_BD7A 812
`define FP16_TO_INDEX_BD78 813
`define FP16_TO_INDEX_BD76 814
`define FP16_TO_INDEX_BD74 815
`define FP16_TO_INDEX_BD72 816
`define FP16_TO_INDEX_BD70 817
`define FP16_TO_INDEX_BD6D 818
`define FP16_TO_INDEX_BD6B 819
`define FP16_TO_INDEX_BD69 820
`define FP16_TO_INDEX_BD67 821
`define FP16_TO_INDEX_BD65 822
`define FP16_TO_INDEX_BD63 823
`define FP16_TO_INDEX_BD61 824
`define FP16_TO_INDEX_BD5F 825
`define FP16_TO_INDEX_BD5D 826
`define FP16_TO_INDEX_BD5B 827
`define FP16_TO_INDEX_BD59 828
`define FP16_TO_INDEX_BD57 829
`define FP16_TO_INDEX_BD55 830
`define FP16_TO_INDEX_BD53 831
`define FP16_TO_INDEX_BD51 832
`define FP16_TO_INDEX_BD4F 833
`define FP16_TO_INDEX_BD4D 834
`define FP16_TO_INDEX_BD4A 835
`define FP16_TO_INDEX_BD48 836
`define FP16_TO_INDEX_BD46 837
`define FP16_TO_INDEX_BD44 838
`define FP16_TO_INDEX_BD42 839
`define FP16_TO_INDEX_BD40 840
`define FP16_TO_INDEX_BD3E 841
`define FP16_TO_INDEX_BD3C 842
`define FP16_TO_INDEX_BD3A 843
`define FP16_TO_INDEX_BD38 844
`define FP16_TO_INDEX_BD36 845
`define FP16_TO_INDEX_BD34 846
`define FP16_TO_INDEX_BD32 847
`define FP16_TO_INDEX_BD30 848
`define FP16_TO_INDEX_BD2E 849
`define FP16_TO_INDEX_BD2C 850
`define FP16_TO_INDEX_BD2A 851
`define FP16_TO_INDEX_BD28 852
`define FP16_TO_INDEX_BD25 853
`define FP16_TO_INDEX_BD23 854
`define FP16_TO_INDEX_BD21 855
`define FP16_TO_INDEX_BD1F 856
`define FP16_TO_INDEX_BD1D 857
`define FP16_TO_INDEX_BD1B 858
`define FP16_TO_INDEX_BD19 859
`define FP16_TO_INDEX_BD17 860
`define FP16_TO_INDEX_BD15 861
`define FP16_TO_INDEX_BD13 862
`define FP16_TO_INDEX_BD11 863
`define FP16_TO_INDEX_BD0F 864
`define FP16_TO_INDEX_BD0D 865
`define FP16_TO_INDEX_BD0B 866
`define FP16_TO_INDEX_BD09 867
`define FP16_TO_INDEX_BD07 868
`define FP16_TO_INDEX_BD05 869
`define FP16_TO_INDEX_BD02 870
`define FP16_TO_INDEX_BD00 871
`define FP16_TO_INDEX_BCFE 872
`define FP16_TO_INDEX_BCFC 873
`define FP16_TO_INDEX_BCFA 874
`define FP16_TO_INDEX_BCF8 875
`define FP16_TO_INDEX_BCF6 876
`define FP16_TO_INDEX_BCF4 877
`define FP16_TO_INDEX_BCF2 878
`define FP16_TO_INDEX_BCF0 879
`define FP16_TO_INDEX_BCEE 880
`define FP16_TO_INDEX_BCEC 881
`define FP16_TO_INDEX_BCEA 882
`define FP16_TO_INDEX_BCE8 883
`define FP16_TO_INDEX_BCE6 884
`define FP16_TO_INDEX_BCE4 885
`define FP16_TO_INDEX_BCE2 886
`define FP16_TO_INDEX_BCE0 887
`define FP16_TO_INDEX_BCDD 888
`define FP16_TO_INDEX_BCDB 889
`define FP16_TO_INDEX_BCD9 890
`define FP16_TO_INDEX_BCD7 891
`define FP16_TO_INDEX_BCD5 892
`define FP16_TO_INDEX_BCD3 893
`define FP16_TO_INDEX_BCD1 894
`define FP16_TO_INDEX_BCCF 895
`define FP16_TO_INDEX_BCCD 896
`define FP16_TO_INDEX_BCCB 897
`define FP16_TO_INDEX_BCC9 898
`define FP16_TO_INDEX_BCC7 899
`define FP16_TO_INDEX_BCC5 900
`define FP16_TO_INDEX_BCC3 901
`define FP16_TO_INDEX_BCC1 902
`define FP16_TO_INDEX_BCBF 903
`define FP16_TO_INDEX_BCBD 904
`define FP16_TO_INDEX_BCBA 905
`define FP16_TO_INDEX_BCB8 906
`define FP16_TO_INDEX_BCB6 907
`define FP16_TO_INDEX_BCB4 908
`define FP16_TO_INDEX_BCB2 909
`define FP16_TO_INDEX_BCB0 910
`define FP16_TO_INDEX_BCAE 911
`define FP16_TO_INDEX_BCAC 912
`define FP16_TO_INDEX_BCAA 913
`define FP16_TO_INDEX_BCA8 914
`define FP16_TO_INDEX_BCA6 915
`define FP16_TO_INDEX_BCA4 916
`define FP16_TO_INDEX_BCA2 917
`define FP16_TO_INDEX_BCA0 918
`define FP16_TO_INDEX_BC9E 919
`define FP16_TO_INDEX_BC9C 920
`define FP16_TO_INDEX_BC9A 921
`define FP16_TO_INDEX_BC98 922
`define FP16_TO_INDEX_BC95 923
`define FP16_TO_INDEX_BC93 924
`define FP16_TO_INDEX_BC91 925
`define FP16_TO_INDEX_BC8F 926
`define FP16_TO_INDEX_BC8D 927
`define FP16_TO_INDEX_BC8B 928
`define FP16_TO_INDEX_BC89 929
`define FP16_TO_INDEX_BC87 930
`define FP16_TO_INDEX_BC85 931
`define FP16_TO_INDEX_BC83 932
`define FP16_TO_INDEX_BC81 933
`define FP16_TO_INDEX_BC7F 934
`define FP16_TO_INDEX_BC7D 935
`define FP16_TO_INDEX_BC7B 936
`define FP16_TO_INDEX_BC79 937
`define FP16_TO_INDEX_BC77 938
`define FP16_TO_INDEX_BC75 939
`define FP16_TO_INDEX_BC73 940
`define FP16_TO_INDEX_BC70 941
`define FP16_TO_INDEX_BC6E 942
`define FP16_TO_INDEX_BC6C 943
`define FP16_TO_INDEX_BC6A 944
`define FP16_TO_INDEX_BC68 945
`define FP16_TO_INDEX_BC66 946
`define FP16_TO_INDEX_BC64 947
`define FP16_TO_INDEX_BC62 948
`define FP16_TO_INDEX_BC60 949
`define FP16_TO_INDEX_BC5E 950
`define FP16_TO_INDEX_BC5C 951
`define FP16_TO_INDEX_BC5A 952
`define FP16_TO_INDEX_BC58 953
`define FP16_TO_INDEX_BC56 954
`define FP16_TO_INDEX_BC54 955
`define FP16_TO_INDEX_BC52 956
`define FP16_TO_INDEX_BC50 957
`define FP16_TO_INDEX_BC4D 958
`define FP16_TO_INDEX_BC4B 959
`define FP16_TO_INDEX_BC49 960
`define FP16_TO_INDEX_BC47 961
`define FP16_TO_INDEX_BC45 962
`define FP16_TO_INDEX_BC43 963
`define FP16_TO_INDEX_BC41 964
`define FP16_TO_INDEX_BC3F 965
`define FP16_TO_INDEX_BC3D 966
`define FP16_TO_INDEX_BC3B 967
`define FP16_TO_INDEX_BC39 968
`define FP16_TO_INDEX_BC37 969
`define FP16_TO_INDEX_BC35 970
`define FP16_TO_INDEX_BC33 971
`define FP16_TO_INDEX_BC31 972
`define FP16_TO_INDEX_BC2F 973
`define FP16_TO_INDEX_BC2D 974
`define FP16_TO_INDEX_BC2B 975
`define FP16_TO_INDEX_BC28 976
`define FP16_TO_INDEX_BC26 977
`define FP16_TO_INDEX_BC24 978
`define FP16_TO_INDEX_BC22 979
`define FP16_TO_INDEX_BC20 980
`define FP16_TO_INDEX_BC1E 981
`define FP16_TO_INDEX_BC1C 982
`define FP16_TO_INDEX_BC1A 983
`define FP16_TO_INDEX_BC18 984
`define FP16_TO_INDEX_BC16 985
`define FP16_TO_INDEX_BC14 986
`define FP16_TO_INDEX_BC12 987
`define FP16_TO_INDEX_BC10 988
`define FP16_TO_INDEX_BC0E 989
`define FP16_TO_INDEX_BC0C 990
`define FP16_TO_INDEX_BC0A 991
`define FP16_TO_INDEX_BC08 992
`define FP16_TO_INDEX_BC05 993
`define FP16_TO_INDEX_BC03 994
`define FP16_TO_INDEX_BC01 995
`define FP16_TO_INDEX_BBFF 996
`define FP16_TO_INDEX_BBFB 997
`define FP16_TO_INDEX_BBF6 998
`define FP16_TO_INDEX_BBF2 999
`define FP16_TO_INDEX_BBEE 1000
`define FP16_TO_INDEX_BBEA 1001
`define FP16_TO_INDEX_BBE6 1002
`define FP16_TO_INDEX_BBE2 1003
`define FP16_TO_INDEX_BBDE 1004
`define FP16_TO_INDEX_BBDA 1005
`define FP16_TO_INDEX_BBD5 1006
`define FP16_TO_INDEX_BBD1 1007
`define FP16_TO_INDEX_BBCD 1008
`define FP16_TO_INDEX_BBC9 1009
`define FP16_TO_INDEX_BBC5 1010
`define FP16_TO_INDEX_BBC1 1011
`define FP16_TO_INDEX_BBBD 1012
`define FP16_TO_INDEX_BBB9 1013
`define FP16_TO_INDEX_BBB5 1014
`define FP16_TO_INDEX_BBB0 1015
`define FP16_TO_INDEX_BBAC 1016
`define FP16_TO_INDEX_BBA8 1017
`define FP16_TO_INDEX_BBA4 1018
`define FP16_TO_INDEX_BBA0 1019
`define FP16_TO_INDEX_BB9C 1020
`define FP16_TO_INDEX_BB98 1021
`define FP16_TO_INDEX_BB94 1022
`define FP16_TO_INDEX_BB90 1023
`define FP16_TO_INDEX_BB8B 1024
`define FP16_TO_INDEX_BB87 1025
`define FP16_TO_INDEX_BB83 1026
`define FP16_TO_INDEX_BB7F 1027
`define FP16_TO_INDEX_BB7B 1028
`define FP16_TO_INDEX_BB77 1029
`define FP16_TO_INDEX_BB73 1030
`define FP16_TO_INDEX_BB6F 1031
`define FP16_TO_INDEX_BB6B 1032
`define FP16_TO_INDEX_BB66 1033
`define FP16_TO_INDEX_BB62 1034
`define FP16_TO_INDEX_BB5E 1035
`define FP16_TO_INDEX_BB5A 1036
`define FP16_TO_INDEX_BB56 1037
`define FP16_TO_INDEX_BB52 1038
`define FP16_TO_INDEX_BB4E 1039
`define FP16_TO_INDEX_BB4A 1040
`define FP16_TO_INDEX_BB46 1041
`define FP16_TO_INDEX_BB41 1042
`define FP16_TO_INDEX_BB3D 1043
`define FP16_TO_INDEX_BB39 1044
`define FP16_TO_INDEX_BB35 1045
`define FP16_TO_INDEX_BB31 1046
`define FP16_TO_INDEX_BB2D 1047
`define FP16_TO_INDEX_BB29 1048
`define FP16_TO_INDEX_BB25 1049
`define FP16_TO_INDEX_BB20 1050
`define FP16_TO_INDEX_BB1C 1051
`define FP16_TO_INDEX_BB18 1052
`define FP16_TO_INDEX_BB14 1053
`define FP16_TO_INDEX_BB10 1054
`define FP16_TO_INDEX_BB0C 1055
`define FP16_TO_INDEX_BB08 1056
`define FP16_TO_INDEX_BB04 1057
`define FP16_TO_INDEX_BB00 1058
`define FP16_TO_INDEX_BAFB 1059
`define FP16_TO_INDEX_BAF7 1060
`define FP16_TO_INDEX_BAF3 1061
`define FP16_TO_INDEX_BAEF 1062
`define FP16_TO_INDEX_BAEB 1063
`define FP16_TO_INDEX_BAE7 1064
`define FP16_TO_INDEX_BAE3 1065
`define FP16_TO_INDEX_BADF 1066
`define FP16_TO_INDEX_BADB 1067
`define FP16_TO_INDEX_BAD6 1068
`define FP16_TO_INDEX_BAD2 1069
`define FP16_TO_INDEX_BACE 1070
`define FP16_TO_INDEX_BACA 1071
`define FP16_TO_INDEX_BAC6 1072
`define FP16_TO_INDEX_BAC2 1073
`define FP16_TO_INDEX_BABE 1074
`define FP16_TO_INDEX_BABA 1075
`define FP16_TO_INDEX_BAB6 1076
`define FP16_TO_INDEX_BAB1 1077
`define FP16_TO_INDEX_BAAD 1078
`define FP16_TO_INDEX_BAA9 1079
`define FP16_TO_INDEX_BAA5 1080
`define FP16_TO_INDEX_BAA1 1081
`define FP16_TO_INDEX_BA9D 1082
`define FP16_TO_INDEX_BA99 1083
`define FP16_TO_INDEX_BA95 1084
`define FP16_TO_INDEX_BA90 1085
`define FP16_TO_INDEX_BA8C 1086
`define FP16_TO_INDEX_BA88 1087
`define FP16_TO_INDEX_BA84 1088
`define FP16_TO_INDEX_BA80 1089
`define FP16_TO_INDEX_BA7C 1090
`define FP16_TO_INDEX_BA78 1091
`define FP16_TO_INDEX_BA74 1092
`define FP16_TO_INDEX_BA70 1093
`define FP16_TO_INDEX_BA6B 1094
`define FP16_TO_INDEX_BA67 1095
`define FP16_TO_INDEX_BA63 1096
`define FP16_TO_INDEX_BA5F 1097
`define FP16_TO_INDEX_BA5B 1098
`define FP16_TO_INDEX_BA57 1099
`define FP16_TO_INDEX_BA53 1100
`define FP16_TO_INDEX_BA4F 1101
`define FP16_TO_INDEX_BA4B 1102
`define FP16_TO_INDEX_BA46 1103
`define FP16_TO_INDEX_BA42 1104
`define FP16_TO_INDEX_BA3E 1105
`define FP16_TO_INDEX_BA3A 1106
`define FP16_TO_INDEX_BA36 1107
`define FP16_TO_INDEX_BA32 1108
`define FP16_TO_INDEX_BA2E 1109
`define FP16_TO_INDEX_BA2A 1110
`define FP16_TO_INDEX_BA26 1111
`define FP16_TO_INDEX_BA21 1112
`define FP16_TO_INDEX_BA1D 1113
`define FP16_TO_INDEX_BA19 1114
`define FP16_TO_INDEX_BA15 1115
`define FP16_TO_INDEX_BA11 1116
`define FP16_TO_INDEX_BA0D 1117
`define FP16_TO_INDEX_BA09 1118
`define FP16_TO_INDEX_BA05 1119
`define FP16_TO_INDEX_BA01 1120
`define FP16_TO_INDEX_B9FC 1121
`define FP16_TO_INDEX_B9F8 1122
`define FP16_TO_INDEX_B9F4 1123
`define FP16_TO_INDEX_B9F0 1124
`define FP16_TO_INDEX_B9EC 1125
`define FP16_TO_INDEX_B9E8 1126
`define FP16_TO_INDEX_B9E4 1127
`define FP16_TO_INDEX_B9E0 1128
`define FP16_TO_INDEX_B9DB 1129
`define FP16_TO_INDEX_B9D7 1130
`define FP16_TO_INDEX_B9D3 1131
`define FP16_TO_INDEX_B9CF 1132
`define FP16_TO_INDEX_B9CB 1133
`define FP16_TO_INDEX_B9C7 1134
`define FP16_TO_INDEX_B9C3 1135
`define FP16_TO_INDEX_B9BF 1136
`define FP16_TO_INDEX_B9BB 1137
`define FP16_TO_INDEX_B9B6 1138
`define FP16_TO_INDEX_B9B2 1139
`define FP16_TO_INDEX_B9AE 1140
`define FP16_TO_INDEX_B9AA 1141
`define FP16_TO_INDEX_B9A6 1142
`define FP16_TO_INDEX_B9A2 1143
`define FP16_TO_INDEX_B99E 1144
`define FP16_TO_INDEX_B99A 1145
`define FP16_TO_INDEX_B996 1146
`define FP16_TO_INDEX_B991 1147
`define FP16_TO_INDEX_B98D 1148
`define FP16_TO_INDEX_B989 1149
`define FP16_TO_INDEX_B985 1150
`define FP16_TO_INDEX_B981 1151
`define FP16_TO_INDEX_B97D 1152
`define FP16_TO_INDEX_B979 1153
`define FP16_TO_INDEX_B975 1154
`define FP16_TO_INDEX_B971 1155
`define FP16_TO_INDEX_B96C 1156
`define FP16_TO_INDEX_B968 1157
`define FP16_TO_INDEX_B964 1158
`define FP16_TO_INDEX_B960 1159
`define FP16_TO_INDEX_B95C 1160
`define FP16_TO_INDEX_B958 1161
`define FP16_TO_INDEX_B954 1162
`define FP16_TO_INDEX_B950 1163
`define FP16_TO_INDEX_B94C 1164
`define FP16_TO_INDEX_B947 1165
`define FP16_TO_INDEX_B943 1166
`define FP16_TO_INDEX_B93F 1167
`define FP16_TO_INDEX_B93B 1168
`define FP16_TO_INDEX_B937 1169
`define FP16_TO_INDEX_B933 1170
`define FP16_TO_INDEX_B92F 1171
`define FP16_TO_INDEX_B92B 1172
`define FP16_TO_INDEX_B926 1173
`define FP16_TO_INDEX_B922 1174
`define FP16_TO_INDEX_B91E 1175
`define FP16_TO_INDEX_B91A 1176
`define FP16_TO_INDEX_B916 1177
`define FP16_TO_INDEX_B912 1178
`define FP16_TO_INDEX_B90E 1179
`define FP16_TO_INDEX_B90A 1180
`define FP16_TO_INDEX_B906 1181
`define FP16_TO_INDEX_B901 1182
`define FP16_TO_INDEX_B8FD 1183
`define FP16_TO_INDEX_B8F9 1184
`define FP16_TO_INDEX_B8F5 1185
`define FP16_TO_INDEX_B8F1 1186
`define FP16_TO_INDEX_B8ED 1187
`define FP16_TO_INDEX_B8E9 1188
`define FP16_TO_INDEX_B8E5 1189
`define FP16_TO_INDEX_B8E1 1190
`define FP16_TO_INDEX_B8DC 1191
`define FP16_TO_INDEX_B8D8 1192
`define FP16_TO_INDEX_B8D4 1193
`define FP16_TO_INDEX_B8D0 1194
`define FP16_TO_INDEX_B8CC 1195
`define FP16_TO_INDEX_B8C8 1196
`define FP16_TO_INDEX_B8C4 1197
`define FP16_TO_INDEX_B8C0 1198
`define FP16_TO_INDEX_B8BC 1199
`define FP16_TO_INDEX_B8B7 1200
`define FP16_TO_INDEX_B8B3 1201
`define FP16_TO_INDEX_B8AF 1202
`define FP16_TO_INDEX_B8AB 1203
`define FP16_TO_INDEX_B8A7 1204
`define FP16_TO_INDEX_B8A3 1205
`define FP16_TO_INDEX_B89F 1206
`define FP16_TO_INDEX_B89B 1207
`define FP16_TO_INDEX_B896 1208
`define FP16_TO_INDEX_B892 1209
`define FP16_TO_INDEX_B88E 1210
`define FP16_TO_INDEX_B88A 1211
`define FP16_TO_INDEX_B886 1212
`define FP16_TO_INDEX_B882 1213
`define FP16_TO_INDEX_B87E 1214
`define FP16_TO_INDEX_B87A 1215
`define FP16_TO_INDEX_B876 1216
`define FP16_TO_INDEX_B871 1217
`define FP16_TO_INDEX_B86D 1218
`define FP16_TO_INDEX_B869 1219
`define FP16_TO_INDEX_B865 1220
`define FP16_TO_INDEX_B861 1221
`define FP16_TO_INDEX_B85D 1222
`define FP16_TO_INDEX_B859 1223
`define FP16_TO_INDEX_B855 1224
`define FP16_TO_INDEX_B851 1225
`define FP16_TO_INDEX_B84C 1226
`define FP16_TO_INDEX_B848 1227
`define FP16_TO_INDEX_B844 1228
`define FP16_TO_INDEX_B840 1229
`define FP16_TO_INDEX_B83C 1230
`define FP16_TO_INDEX_B838 1231
`define FP16_TO_INDEX_B834 1232
`define FP16_TO_INDEX_B830 1233
`define FP16_TO_INDEX_B82C 1234
`define FP16_TO_INDEX_B827 1235
`define FP16_TO_INDEX_B823 1236
`define FP16_TO_INDEX_B81F 1237
`define FP16_TO_INDEX_B81B 1238
`define FP16_TO_INDEX_B817 1239
`define FP16_TO_INDEX_B813 1240
`define FP16_TO_INDEX_B80F 1241
`define FP16_TO_INDEX_B80B 1242
`define FP16_TO_INDEX_B807 1243
`define FP16_TO_INDEX_B802 1244
`define FP16_TO_INDEX_B7FD 1245
`define FP16_TO_INDEX_B7F4 1246
`define FP16_TO_INDEX_B7EC 1247
`define FP16_TO_INDEX_B7E4 1248
`define FP16_TO_INDEX_B7DC 1249
`define FP16_TO_INDEX_B7D3 1250
`define FP16_TO_INDEX_B7CB 1251
`define FP16_TO_INDEX_B7C3 1252
`define FP16_TO_INDEX_B7BB 1253
`define FP16_TO_INDEX_B7B3 1254
`define FP16_TO_INDEX_B7AA 1255
`define FP16_TO_INDEX_B7A2 1256
`define FP16_TO_INDEX_B79A 1257
`define FP16_TO_INDEX_B792 1258
`define FP16_TO_INDEX_B789 1259
`define FP16_TO_INDEX_B781 1260
`define FP16_TO_INDEX_B779 1261
`define FP16_TO_INDEX_B771 1262
`define FP16_TO_INDEX_B768 1263
`define FP16_TO_INDEX_B760 1264
`define FP16_TO_INDEX_B758 1265
`define FP16_TO_INDEX_B750 1266
`define FP16_TO_INDEX_B748 1267
`define FP16_TO_INDEX_B73F 1268
`define FP16_TO_INDEX_B737 1269
`define FP16_TO_INDEX_B72F 1270
`define FP16_TO_INDEX_B727 1271
`define FP16_TO_INDEX_B71E 1272
`define FP16_TO_INDEX_B716 1273
`define FP16_TO_INDEX_B70E 1274
`define FP16_TO_INDEX_B706 1275
`define FP16_TO_INDEX_B6FE 1276
`define FP16_TO_INDEX_B6F5 1277
`define FP16_TO_INDEX_B6ED 1278
`define FP16_TO_INDEX_B6E5 1279
`define FP16_TO_INDEX_B6DD 1280
`define FP16_TO_INDEX_B6D4 1281
`define FP16_TO_INDEX_B6CC 1282
`define FP16_TO_INDEX_B6C4 1283
`define FP16_TO_INDEX_B6BC 1284
`define FP16_TO_INDEX_B6B3 1285
`define FP16_TO_INDEX_B6AB 1286
`define FP16_TO_INDEX_B6A3 1287
`define FP16_TO_INDEX_B69B 1288
`define FP16_TO_INDEX_B693 1289
`define FP16_TO_INDEX_B68A 1290
`define FP16_TO_INDEX_B682 1291
`define FP16_TO_INDEX_B67A 1292
`define FP16_TO_INDEX_B672 1293
`define FP16_TO_INDEX_B669 1294
`define FP16_TO_INDEX_B661 1295
`define FP16_TO_INDEX_B659 1296
`define FP16_TO_INDEX_B651 1297
`define FP16_TO_INDEX_B649 1298
`define FP16_TO_INDEX_B640 1299
`define FP16_TO_INDEX_B638 1300
`define FP16_TO_INDEX_B630 1301
`define FP16_TO_INDEX_B628 1302
`define FP16_TO_INDEX_B61F 1303
`define FP16_TO_INDEX_B617 1304
`define FP16_TO_INDEX_B60F 1305
`define FP16_TO_INDEX_B607 1306
`define FP16_TO_INDEX_B5FE 1307
`define FP16_TO_INDEX_B5F6 1308
`define FP16_TO_INDEX_B5EE 1309
`define FP16_TO_INDEX_B5E6 1310
`define FP16_TO_INDEX_B5DE 1311
`define FP16_TO_INDEX_B5D5 1312
`define FP16_TO_INDEX_B5CD 1313
`define FP16_TO_INDEX_B5C5 1314
`define FP16_TO_INDEX_B5BD 1315
`define FP16_TO_INDEX_B5B4 1316
`define FP16_TO_INDEX_B5AC 1317
`define FP16_TO_INDEX_B5A4 1318
`define FP16_TO_INDEX_B59C 1319
`define FP16_TO_INDEX_B593 1320
`define FP16_TO_INDEX_B58B 1321
`define FP16_TO_INDEX_B583 1322
`define FP16_TO_INDEX_B57B 1323
`define FP16_TO_INDEX_B573 1324
`define FP16_TO_INDEX_B56A 1325
`define FP16_TO_INDEX_B562 1326
`define FP16_TO_INDEX_B55A 1327
`define FP16_TO_INDEX_B552 1328
`define FP16_TO_INDEX_B549 1329
`define FP16_TO_INDEX_B541 1330
`define FP16_TO_INDEX_B539 1331
`define FP16_TO_INDEX_B531 1332
`define FP16_TO_INDEX_B529 1333
`define FP16_TO_INDEX_B520 1334
`define FP16_TO_INDEX_B518 1335
`define FP16_TO_INDEX_B510 1336
`define FP16_TO_INDEX_B508 1337
`define FP16_TO_INDEX_B4FF 1338
`define FP16_TO_INDEX_B4F7 1339
`define FP16_TO_INDEX_B4EF 1340
`define FP16_TO_INDEX_B4E7 1341
`define FP16_TO_INDEX_B4DE 1342
`define FP16_TO_INDEX_B4D6 1343
`define FP16_TO_INDEX_B4CE 1344
`define FP16_TO_INDEX_B4C6 1345
`define FP16_TO_INDEX_B4BE 1346
`define FP16_TO_INDEX_B4B5 1347
`define FP16_TO_INDEX_B4AD 1348
`define FP16_TO_INDEX_B4A5 1349
`define FP16_TO_INDEX_B49D 1350
`define FP16_TO_INDEX_B494 1351
`define FP16_TO_INDEX_B48C 1352
`define FP16_TO_INDEX_B484 1353
`define FP16_TO_INDEX_B47C 1354
`define FP16_TO_INDEX_B474 1355
`define FP16_TO_INDEX_B46B 1356
`define FP16_TO_INDEX_B463 1357
`define FP16_TO_INDEX_B45B 1358
`define FP16_TO_INDEX_B453 1359
`define FP16_TO_INDEX_B44A 1360
`define FP16_TO_INDEX_B442 1361
`define FP16_TO_INDEX_B43A 1362
`define FP16_TO_INDEX_B432 1363
`define FP16_TO_INDEX_B429 1364
`define FP16_TO_INDEX_B421 1365
`define FP16_TO_INDEX_B419 1366
`define FP16_TO_INDEX_B411 1367
`define FP16_TO_INDEX_B409 1368
`define FP16_TO_INDEX_B400 1369
`define FP16_TO_INDEX_B3F0 1370
`define FP16_TO_INDEX_B3E0 1371
`define FP16_TO_INDEX_B3CF 1372
`define FP16_TO_INDEX_B3BF 1373
`define FP16_TO_INDEX_B3AE 1374
`define FP16_TO_INDEX_B39E 1375
`define FP16_TO_INDEX_B38D 1376
`define FP16_TO_INDEX_B37D 1377
`define FP16_TO_INDEX_B36D 1378
`define FP16_TO_INDEX_B35C 1379
`define FP16_TO_INDEX_B34C 1380
`define FP16_TO_INDEX_B33B 1381
`define FP16_TO_INDEX_B32B 1382
`define FP16_TO_INDEX_B31A 1383
`define FP16_TO_INDEX_B30A 1384
`define FP16_TO_INDEX_B2F9 1385
`define FP16_TO_INDEX_B2E9 1386
`define FP16_TO_INDEX_B2D8 1387
`define FP16_TO_INDEX_B2C8 1388
`define FP16_TO_INDEX_B2B8 1389
`define FP16_TO_INDEX_B2A7 1390
`define FP16_TO_INDEX_B297 1391
`define FP16_TO_INDEX_B286 1392
`define FP16_TO_INDEX_B276 1393
`define FP16_TO_INDEX_B265 1394
`define FP16_TO_INDEX_B255 1395
`define FP16_TO_INDEX_B244 1396
`define FP16_TO_INDEX_B234 1397
`define FP16_TO_INDEX_B223 1398
`define FP16_TO_INDEX_B213 1399
`define FP16_TO_INDEX_B203 1400
`define FP16_TO_INDEX_B1F2 1401
`define FP16_TO_INDEX_B1E2 1402
`define FP16_TO_INDEX_B1D1 1403
`define FP16_TO_INDEX_B1C1 1404
`define FP16_TO_INDEX_B1B0 1405
`define FP16_TO_INDEX_B1A0 1406
`define FP16_TO_INDEX_B18F 1407
`define FP16_TO_INDEX_B17F 1408
`define FP16_TO_INDEX_B16E 1409
`define FP16_TO_INDEX_B15E 1410
`define FP16_TO_INDEX_B14E 1411
`define FP16_TO_INDEX_B13D 1412
`define FP16_TO_INDEX_B12D 1413
`define FP16_TO_INDEX_B11C 1414
`define FP16_TO_INDEX_B10C 1415
`define FP16_TO_INDEX_B0FB 1416
`define FP16_TO_INDEX_B0EB 1417
`define FP16_TO_INDEX_B0DA 1418
`define FP16_TO_INDEX_B0CA 1419
`define FP16_TO_INDEX_B0B9 1420
`define FP16_TO_INDEX_B0A9 1421
`define FP16_TO_INDEX_B099 1422
`define FP16_TO_INDEX_B088 1423
`define FP16_TO_INDEX_B078 1424
`define FP16_TO_INDEX_B067 1425
`define FP16_TO_INDEX_B057 1426
`define FP16_TO_INDEX_B046 1427
`define FP16_TO_INDEX_B036 1428
`define FP16_TO_INDEX_B025 1429
`define FP16_TO_INDEX_B015 1430
`define FP16_TO_INDEX_B004 1431
`define FP16_TO_INDEX_AFE8 1432
`define FP16_TO_INDEX_AFC7 1433
`define FP16_TO_INDEX_AFA6 1434
`define FP16_TO_INDEX_AF85 1435
`define FP16_TO_INDEX_AF64 1436
`define FP16_TO_INDEX_AF43 1437
`define FP16_TO_INDEX_AF23 1438
`define FP16_TO_INDEX_AF02 1439
`define FP16_TO_INDEX_AEE1 1440
`define FP16_TO_INDEX_AEC0 1441
`define FP16_TO_INDEX_AE9F 1442
`define FP16_TO_INDEX_AE7E 1443
`define FP16_TO_INDEX_AE5D 1444
`define FP16_TO_INDEX_AE3C 1445
`define FP16_TO_INDEX_AE1B 1446
`define FP16_TO_INDEX_ADFA 1447
`define FP16_TO_INDEX_ADD9 1448
`define FP16_TO_INDEX_ADB9 1449
`define FP16_TO_INDEX_AD98 1450
`define FP16_TO_INDEX_AD77 1451
`define FP16_TO_INDEX_AD56 1452
`define FP16_TO_INDEX_AD35 1453
`define FP16_TO_INDEX_AD14 1454
`define FP16_TO_INDEX_ACF3 1455
`define FP16_TO_INDEX_ACD2 1456
`define FP16_TO_INDEX_ACB1 1457
`define FP16_TO_INDEX_AC90 1458
`define FP16_TO_INDEX_AC6F 1459
`define FP16_TO_INDEX_AC4F 1460
`define FP16_TO_INDEX_AC2E 1461
`define FP16_TO_INDEX_AC0D 1462
`define FP16_TO_INDEX_ABD8 1463
`define FP16_TO_INDEX_AB96 1464
`define FP16_TO_INDEX_AB54 1465
`define FP16_TO_INDEX_AB12 1466
`define FP16_TO_INDEX_AAD0 1467
`define FP16_TO_INDEX_AA8E 1468
`define FP16_TO_INDEX_AA4D 1469
`define FP16_TO_INDEX_AA0B 1470
`define FP16_TO_INDEX_A9C9 1471
`define FP16_TO_INDEX_A987 1472
`define FP16_TO_INDEX_A945 1473
`define FP16_TO_INDEX_A904 1474
`define FP16_TO_INDEX_A8C2 1475
`define FP16_TO_INDEX_A880 1476
`define FP16_TO_INDEX_A83E 1477
`define FP16_TO_INDEX_A7F8 1478
`define FP16_TO_INDEX_A775 1479
`define FP16_TO_INDEX_A6F1 1480
`define FP16_TO_INDEX_A66E 1481
`define FP16_TO_INDEX_A5EA 1482
`define FP16_TO_INDEX_A566 1483
`define FP16_TO_INDEX_A4E3 1484
`define FP16_TO_INDEX_A45F 1485
`define FP16_TO_INDEX_A3B7 1486
`define FP16_TO_INDEX_A2AF 1487
`define FP16_TO_INDEX_A1A8 1488
`define FP16_TO_INDEX_A0A1 1489
`define FP16_TO_INDEX_9F33 1490
`define FP16_TO_INDEX_9D24 1491
`define FP16_TO_INDEX_9A2C 1492
`define FP16_TO_INDEX_941D 1493
`define FP16_TO_INDEX_141D 1494
`define FP16_TO_INDEX_1A2C 1495
`define FP16_TO_INDEX_1D24 1496
`define FP16_TO_INDEX_1F33 1497
`define FP16_TO_INDEX_20A1 1498
`define FP16_TO_INDEX_21A8 1499
`define FP16_TO_INDEX_22AF 1500
`define FP16_TO_INDEX_23B7 1501
`define FP16_TO_INDEX_245F 1502
`define FP16_TO_INDEX_24E3 1503
`define FP16_TO_INDEX_2566 1504
`define FP16_TO_INDEX_25EA 1505
`define FP16_TO_INDEX_266E 1506
`define FP16_TO_INDEX_26F1 1507
`define FP16_TO_INDEX_2775 1508
`define FP16_TO_INDEX_27F8 1509
`define FP16_TO_INDEX_283E 1510
`define FP16_TO_INDEX_2880 1511
`define FP16_TO_INDEX_28C2 1512
`define FP16_TO_INDEX_2904 1513
`define FP16_TO_INDEX_2945 1514
`define FP16_TO_INDEX_2987 1515
`define FP16_TO_INDEX_29C9 1516
`define FP16_TO_INDEX_2A0B 1517
`define FP16_TO_INDEX_2A4D 1518
`define FP16_TO_INDEX_2A8E 1519
`define FP16_TO_INDEX_2AD0 1520
`define FP16_TO_INDEX_2B12 1521
`define FP16_TO_INDEX_2B54 1522
`define FP16_TO_INDEX_2B96 1523
`define FP16_TO_INDEX_2BD8 1524
`define FP16_TO_INDEX_2C0D 1525
`define FP16_TO_INDEX_2C2E 1526
`define FP16_TO_INDEX_2C4F 1527
`define FP16_TO_INDEX_2C6F 1528
`define FP16_TO_INDEX_2C90 1529
`define FP16_TO_INDEX_2CB1 1530
`define FP16_TO_INDEX_2CD2 1531
`define FP16_TO_INDEX_2CF3 1532
`define FP16_TO_INDEX_2D14 1533
`define FP16_TO_INDEX_2D35 1534
`define FP16_TO_INDEX_2D56 1535
`define FP16_TO_INDEX_2D77 1536
`define FP16_TO_INDEX_2D98 1537
`define FP16_TO_INDEX_2DB9 1538
`define FP16_TO_INDEX_2DD9 1539
`define FP16_TO_INDEX_2DFA 1540
`define FP16_TO_INDEX_2E1B 1541
`define FP16_TO_INDEX_2E3C 1542
`define FP16_TO_INDEX_2E5D 1543
`define FP16_TO_INDEX_2E7E 1544
`define FP16_TO_INDEX_2E9F 1545
`define FP16_TO_INDEX_2EC0 1546
`define FP16_TO_INDEX_2EE1 1547
`define FP16_TO_INDEX_2F02 1548
`define FP16_TO_INDEX_2F23 1549
`define FP16_TO_INDEX_2F43 1550
`define FP16_TO_INDEX_2F64 1551
`define FP16_TO_INDEX_2F85 1552
`define FP16_TO_INDEX_2FA6 1553
`define FP16_TO_INDEX_2FC7 1554
`define FP16_TO_INDEX_2FE8 1555
`define FP16_TO_INDEX_3004 1556
`define FP16_TO_INDEX_3015 1557
`define FP16_TO_INDEX_3025 1558
`define FP16_TO_INDEX_3036 1559
`define FP16_TO_INDEX_3046 1560
`define FP16_TO_INDEX_3057 1561
`define FP16_TO_INDEX_3067 1562
`define FP16_TO_INDEX_3078 1563
`define FP16_TO_INDEX_3088 1564
`define FP16_TO_INDEX_3099 1565
`define FP16_TO_INDEX_30A9 1566
`define FP16_TO_INDEX_30B9 1567
`define FP16_TO_INDEX_30CA 1568
`define FP16_TO_INDEX_30DA 1569
`define FP16_TO_INDEX_30EB 1570
`define FP16_TO_INDEX_30FB 1571
`define FP16_TO_INDEX_310C 1572
`define FP16_TO_INDEX_311C 1573
`define FP16_TO_INDEX_312D 1574
`define FP16_TO_INDEX_313D 1575
`define FP16_TO_INDEX_314E 1576
`define FP16_TO_INDEX_315E 1577
`define FP16_TO_INDEX_316E 1578
`define FP16_TO_INDEX_317F 1579
`define FP16_TO_INDEX_318F 1580
`define FP16_TO_INDEX_31A0 1581
`define FP16_TO_INDEX_31B0 1582
`define FP16_TO_INDEX_31C1 1583
`define FP16_TO_INDEX_31D1 1584
`define FP16_TO_INDEX_31E2 1585
`define FP16_TO_INDEX_31F2 1586
`define FP16_TO_INDEX_3203 1587
`define FP16_TO_INDEX_3213 1588
`define FP16_TO_INDEX_3223 1589
`define FP16_TO_INDEX_3234 1590
`define FP16_TO_INDEX_3244 1591
`define FP16_TO_INDEX_3255 1592
`define FP16_TO_INDEX_3265 1593
`define FP16_TO_INDEX_3276 1594
`define FP16_TO_INDEX_3286 1595
`define FP16_TO_INDEX_3297 1596
`define FP16_TO_INDEX_32A7 1597
`define FP16_TO_INDEX_32B8 1598
`define FP16_TO_INDEX_32C8 1599
`define FP16_TO_INDEX_32D8 1600
`define FP16_TO_INDEX_32E9 1601
`define FP16_TO_INDEX_32F9 1602
`define FP16_TO_INDEX_330A 1603
`define FP16_TO_INDEX_331A 1604
`define FP16_TO_INDEX_332B 1605
`define FP16_TO_INDEX_333B 1606
`define FP16_TO_INDEX_334C 1607
`define FP16_TO_INDEX_335C 1608
`define FP16_TO_INDEX_336D 1609
`define FP16_TO_INDEX_337D 1610
`define FP16_TO_INDEX_338D 1611
`define FP16_TO_INDEX_339E 1612
`define FP16_TO_INDEX_33AE 1613
`define FP16_TO_INDEX_33BF 1614
`define FP16_TO_INDEX_33CF 1615
`define FP16_TO_INDEX_33E0 1616
`define FP16_TO_INDEX_33F0 1617
`define FP16_TO_INDEX_3400 1618
`define FP16_TO_INDEX_3409 1619
`define FP16_TO_INDEX_3411 1620
`define FP16_TO_INDEX_3419 1621
`define FP16_TO_INDEX_3421 1622
`define FP16_TO_INDEX_3429 1623
`define FP16_TO_INDEX_3432 1624
`define FP16_TO_INDEX_343A 1625
`define FP16_TO_INDEX_3442 1626
`define FP16_TO_INDEX_344A 1627
`define FP16_TO_INDEX_3453 1628
`define FP16_TO_INDEX_345B 1629
`define FP16_TO_INDEX_3463 1630
`define FP16_TO_INDEX_346B 1631
`define FP16_TO_INDEX_3474 1632
`define FP16_TO_INDEX_347C 1633
`define FP16_TO_INDEX_3484 1634
`define FP16_TO_INDEX_348C 1635
`define FP16_TO_INDEX_3494 1636
`define FP16_TO_INDEX_349D 1637
`define FP16_TO_INDEX_34A5 1638
`define FP16_TO_INDEX_34AD 1639
`define FP16_TO_INDEX_34B5 1640
`define FP16_TO_INDEX_34BE 1641
`define FP16_TO_INDEX_34C6 1642
`define FP16_TO_INDEX_34CE 1643
`define FP16_TO_INDEX_34D6 1644
`define FP16_TO_INDEX_34DE 1645
`define FP16_TO_INDEX_34E7 1646
`define FP16_TO_INDEX_34EF 1647
`define FP16_TO_INDEX_34F7 1648
`define FP16_TO_INDEX_34FF 1649
`define FP16_TO_INDEX_3508 1650
`define FP16_TO_INDEX_3510 1651
`define FP16_TO_INDEX_3518 1652
`define FP16_TO_INDEX_3520 1653
`define FP16_TO_INDEX_3529 1654
`define FP16_TO_INDEX_3531 1655
`define FP16_TO_INDEX_3539 1656
`define FP16_TO_INDEX_3541 1657
`define FP16_TO_INDEX_3549 1658
`define FP16_TO_INDEX_3552 1659
`define FP16_TO_INDEX_355A 1660
`define FP16_TO_INDEX_3562 1661
`define FP16_TO_INDEX_356A 1662
`define FP16_TO_INDEX_3573 1663
`define FP16_TO_INDEX_357B 1664
`define FP16_TO_INDEX_3583 1665
`define FP16_TO_INDEX_358B 1666
`define FP16_TO_INDEX_3593 1667
`define FP16_TO_INDEX_359C 1668
`define FP16_TO_INDEX_35A4 1669
`define FP16_TO_INDEX_35AC 1670
`define FP16_TO_INDEX_35B4 1671
`define FP16_TO_INDEX_35BD 1672
`define FP16_TO_INDEX_35C5 1673
`define FP16_TO_INDEX_35CD 1674
`define FP16_TO_INDEX_35D5 1675
`define FP16_TO_INDEX_35DE 1676
`define FP16_TO_INDEX_35E6 1677
`define FP16_TO_INDEX_35EE 1678
`define FP16_TO_INDEX_35F6 1679
`define FP16_TO_INDEX_35FE 1680
`define FP16_TO_INDEX_3607 1681
`define FP16_TO_INDEX_360F 1682
`define FP16_TO_INDEX_3617 1683
`define FP16_TO_INDEX_361F 1684
`define FP16_TO_INDEX_3628 1685
`define FP16_TO_INDEX_3630 1686
`define FP16_TO_INDEX_3638 1687
`define FP16_TO_INDEX_3640 1688
`define FP16_TO_INDEX_3649 1689
`define FP16_TO_INDEX_3651 1690
`define FP16_TO_INDEX_3659 1691
`define FP16_TO_INDEX_3661 1692
`define FP16_TO_INDEX_3669 1693
`define FP16_TO_INDEX_3672 1694
`define FP16_TO_INDEX_367A 1695
`define FP16_TO_INDEX_3682 1696
`define FP16_TO_INDEX_368A 1697
`define FP16_TO_INDEX_3693 1698
`define FP16_TO_INDEX_369B 1699
`define FP16_TO_INDEX_36A3 1700
`define FP16_TO_INDEX_36AB 1701
`define FP16_TO_INDEX_36B3 1702
`define FP16_TO_INDEX_36BC 1703
`define FP16_TO_INDEX_36C4 1704
`define FP16_TO_INDEX_36CC 1705
`define FP16_TO_INDEX_36D4 1706
`define FP16_TO_INDEX_36DD 1707
`define FP16_TO_INDEX_36E5 1708
`define FP16_TO_INDEX_36ED 1709
`define FP16_TO_INDEX_36F5 1710
`define FP16_TO_INDEX_36FE 1711
`define FP16_TO_INDEX_3706 1712
`define FP16_TO_INDEX_370E 1713
`define FP16_TO_INDEX_3716 1714
`define FP16_TO_INDEX_371E 1715
`define FP16_TO_INDEX_3727 1716
`define FP16_TO_INDEX_372F 1717
`define FP16_TO_INDEX_3737 1718
`define FP16_TO_INDEX_373F 1719
`define FP16_TO_INDEX_3748 1720
`define FP16_TO_INDEX_3750 1721
`define FP16_TO_INDEX_3758 1722
`define FP16_TO_INDEX_3760 1723
`define FP16_TO_INDEX_3768 1724
`define FP16_TO_INDEX_3771 1725
`define FP16_TO_INDEX_3779 1726
`define FP16_TO_INDEX_3781 1727
`define FP16_TO_INDEX_3789 1728
`define FP16_TO_INDEX_3792 1729
`define FP16_TO_INDEX_379A 1730
`define FP16_TO_INDEX_37A2 1731
`define FP16_TO_INDEX_37AA 1732
`define FP16_TO_INDEX_37B3 1733
`define FP16_TO_INDEX_37BB 1734
`define FP16_TO_INDEX_37C3 1735
`define FP16_TO_INDEX_37CB 1736
`define FP16_TO_INDEX_37D3 1737
`define FP16_TO_INDEX_37DC 1738
`define FP16_TO_INDEX_37E4 1739
`define FP16_TO_INDEX_37EC 1740
`define FP16_TO_INDEX_37F4 1741
`define FP16_TO_INDEX_37FD 1742
`define FP16_TO_INDEX_3802 1743
`define FP16_TO_INDEX_3807 1744
`define FP16_TO_INDEX_380B 1745
`define FP16_TO_INDEX_380F 1746
`define FP16_TO_INDEX_3813 1747
`define FP16_TO_INDEX_3817 1748
`define FP16_TO_INDEX_381B 1749
`define FP16_TO_INDEX_381F 1750
`define FP16_TO_INDEX_3823 1751
`define FP16_TO_INDEX_3827 1752
`define FP16_TO_INDEX_382C 1753
`define FP16_TO_INDEX_3830 1754
`define FP16_TO_INDEX_3834 1755
`define FP16_TO_INDEX_3838 1756
`define FP16_TO_INDEX_383C 1757
`define FP16_TO_INDEX_3840 1758
`define FP16_TO_INDEX_3844 1759
`define FP16_TO_INDEX_3848 1760
`define FP16_TO_INDEX_384C 1761
`define FP16_TO_INDEX_3851 1762
`define FP16_TO_INDEX_3855 1763
`define FP16_TO_INDEX_3859 1764
`define FP16_TO_INDEX_385D 1765
`define FP16_TO_INDEX_3861 1766
`define FP16_TO_INDEX_3865 1767
`define FP16_TO_INDEX_3869 1768
`define FP16_TO_INDEX_386D 1769
`define FP16_TO_INDEX_3871 1770
`define FP16_TO_INDEX_3876 1771
`define FP16_TO_INDEX_387A 1772
`define FP16_TO_INDEX_387E 1773
`define FP16_TO_INDEX_3882 1774
`define FP16_TO_INDEX_3886 1775
`define FP16_TO_INDEX_388A 1776
`define FP16_TO_INDEX_388E 1777
`define FP16_TO_INDEX_3892 1778
`define FP16_TO_INDEX_3896 1779
`define FP16_TO_INDEX_389B 1780
`define FP16_TO_INDEX_389F 1781
`define FP16_TO_INDEX_38A3 1782
`define FP16_TO_INDEX_38A7 1783
`define FP16_TO_INDEX_38AB 1784
`define FP16_TO_INDEX_38AF 1785
`define FP16_TO_INDEX_38B3 1786
`define FP16_TO_INDEX_38B7 1787
`define FP16_TO_INDEX_38BC 1788
`define FP16_TO_INDEX_38C0 1789
`define FP16_TO_INDEX_38C4 1790
`define FP16_TO_INDEX_38C8 1791
`define FP16_TO_INDEX_38CC 1792
`define FP16_TO_INDEX_38D0 1793
`define FP16_TO_INDEX_38D4 1794
`define FP16_TO_INDEX_38D8 1795
`define FP16_TO_INDEX_38DC 1796
`define FP16_TO_INDEX_38E1 1797
`define FP16_TO_INDEX_38E5 1798
`define FP16_TO_INDEX_38E9 1799
`define FP16_TO_INDEX_38ED 1800
`define FP16_TO_INDEX_38F1 1801
`define FP16_TO_INDEX_38F5 1802
`define FP16_TO_INDEX_38F9 1803
`define FP16_TO_INDEX_38FD 1804
`define FP16_TO_INDEX_3901 1805
`define FP16_TO_INDEX_3906 1806
`define FP16_TO_INDEX_390A 1807
`define FP16_TO_INDEX_390E 1808
`define FP16_TO_INDEX_3912 1809
`define FP16_TO_INDEX_3916 1810
`define FP16_TO_INDEX_391A 1811
`define FP16_TO_INDEX_391E 1812
`define FP16_TO_INDEX_3922 1813
`define FP16_TO_INDEX_3926 1814
`define FP16_TO_INDEX_392B 1815
`define FP16_TO_INDEX_392F 1816
`define FP16_TO_INDEX_3933 1817
`define FP16_TO_INDEX_3937 1818
`define FP16_TO_INDEX_393B 1819
`define FP16_TO_INDEX_393F 1820
`define FP16_TO_INDEX_3943 1821
`define FP16_TO_INDEX_3947 1822
`define FP16_TO_INDEX_394C 1823
`define FP16_TO_INDEX_3950 1824
`define FP16_TO_INDEX_3954 1825
`define FP16_TO_INDEX_3958 1826
`define FP16_TO_INDEX_395C 1827
`define FP16_TO_INDEX_3960 1828
`define FP16_TO_INDEX_3964 1829
`define FP16_TO_INDEX_3968 1830
`define FP16_TO_INDEX_396C 1831
`define FP16_TO_INDEX_3971 1832
`define FP16_TO_INDEX_3975 1833
`define FP16_TO_INDEX_3979 1834
`define FP16_TO_INDEX_397D 1835
`define FP16_TO_INDEX_3981 1836
`define FP16_TO_INDEX_3985 1837
`define FP16_TO_INDEX_3989 1838
`define FP16_TO_INDEX_398D 1839
`define FP16_TO_INDEX_3991 1840
`define FP16_TO_INDEX_3996 1841
`define FP16_TO_INDEX_399A 1842
`define FP16_TO_INDEX_399E 1843
`define FP16_TO_INDEX_39A2 1844
`define FP16_TO_INDEX_39A6 1845
`define FP16_TO_INDEX_39AA 1846
`define FP16_TO_INDEX_39AE 1847
`define FP16_TO_INDEX_39B2 1848
`define FP16_TO_INDEX_39B6 1849
`define FP16_TO_INDEX_39BB 1850
`define FP16_TO_INDEX_39BF 1851
`define FP16_TO_INDEX_39C3 1852
`define FP16_TO_INDEX_39C7 1853
`define FP16_TO_INDEX_39CB 1854
`define FP16_TO_INDEX_39CF 1855
`define FP16_TO_INDEX_39D3 1856
`define FP16_TO_INDEX_39D7 1857
`define FP16_TO_INDEX_39DB 1858
`define FP16_TO_INDEX_39E0 1859
`define FP16_TO_INDEX_39E4 1860
`define FP16_TO_INDEX_39E8 1861
`define FP16_TO_INDEX_39EC 1862
`define FP16_TO_INDEX_39F0 1863
`define FP16_TO_INDEX_39F4 1864
`define FP16_TO_INDEX_39F8 1865
`define FP16_TO_INDEX_39FC 1866
`define FP16_TO_INDEX_3A01 1867
`define FP16_TO_INDEX_3A05 1868
`define FP16_TO_INDEX_3A09 1869
`define FP16_TO_INDEX_3A0D 1870
`define FP16_TO_INDEX_3A11 1871
`define FP16_TO_INDEX_3A15 1872
`define FP16_TO_INDEX_3A19 1873
`define FP16_TO_INDEX_3A1D 1874
`define FP16_TO_INDEX_3A21 1875
`define FP16_TO_INDEX_3A26 1876
`define FP16_TO_INDEX_3A2A 1877
`define FP16_TO_INDEX_3A2E 1878
`define FP16_TO_INDEX_3A32 1879
`define FP16_TO_INDEX_3A36 1880
`define FP16_TO_INDEX_3A3A 1881
`define FP16_TO_INDEX_3A3E 1882
`define FP16_TO_INDEX_3A42 1883
`define FP16_TO_INDEX_3A46 1884
`define FP16_TO_INDEX_3A4B 1885
`define FP16_TO_INDEX_3A4F 1886
`define FP16_TO_INDEX_3A53 1887
`define FP16_TO_INDEX_3A57 1888
`define FP16_TO_INDEX_3A5B 1889
`define FP16_TO_INDEX_3A5F 1890
`define FP16_TO_INDEX_3A63 1891
`define FP16_TO_INDEX_3A67 1892
`define FP16_TO_INDEX_3A6B 1893
`define FP16_TO_INDEX_3A70 1894
`define FP16_TO_INDEX_3A74 1895
`define FP16_TO_INDEX_3A78 1896
`define FP16_TO_INDEX_3A7C 1897
`define FP16_TO_INDEX_3A80 1898
`define FP16_TO_INDEX_3A84 1899
`define FP16_TO_INDEX_3A88 1900
`define FP16_TO_INDEX_3A8C 1901
`define FP16_TO_INDEX_3A90 1902
`define FP16_TO_INDEX_3A95 1903
`define FP16_TO_INDEX_3A99 1904
`define FP16_TO_INDEX_3A9D 1905
`define FP16_TO_INDEX_3AA1 1906
`define FP16_TO_INDEX_3AA5 1907
`define FP16_TO_INDEX_3AA9 1908
`define FP16_TO_INDEX_3AAD 1909
`define FP16_TO_INDEX_3AB1 1910
`define FP16_TO_INDEX_3AB6 1911
`define FP16_TO_INDEX_3ABA 1912
`define FP16_TO_INDEX_3ABE 1913
`define FP16_TO_INDEX_3AC2 1914
`define FP16_TO_INDEX_3AC6 1915
`define FP16_TO_INDEX_3ACA 1916
`define FP16_TO_INDEX_3ACE 1917
`define FP16_TO_INDEX_3AD2 1918
`define FP16_TO_INDEX_3AD6 1919
`define FP16_TO_INDEX_3ADB 1920
`define FP16_TO_INDEX_3ADF 1921
`define FP16_TO_INDEX_3AE3 1922
`define FP16_TO_INDEX_3AE7 1923
`define FP16_TO_INDEX_3AEB 1924
`define FP16_TO_INDEX_3AEF 1925
`define FP16_TO_INDEX_3AF3 1926
`define FP16_TO_INDEX_3AF7 1927
`define FP16_TO_INDEX_3AFB 1928
`define FP16_TO_INDEX_3B00 1929
`define FP16_TO_INDEX_3B04 1930
`define FP16_TO_INDEX_3B08 1931
`define FP16_TO_INDEX_3B0C 1932
`define FP16_TO_INDEX_3B10 1933
`define FP16_TO_INDEX_3B14 1934
`define FP16_TO_INDEX_3B18 1935
`define FP16_TO_INDEX_3B1C 1936
`define FP16_TO_INDEX_3B20 1937
`define FP16_TO_INDEX_3B25 1938
`define FP16_TO_INDEX_3B29 1939
`define FP16_TO_INDEX_3B2D 1940
`define FP16_TO_INDEX_3B31 1941
`define FP16_TO_INDEX_3B35 1942
`define FP16_TO_INDEX_3B39 1943
`define FP16_TO_INDEX_3B3D 1944
`define FP16_TO_INDEX_3B41 1945
`define FP16_TO_INDEX_3B46 1946
`define FP16_TO_INDEX_3B4A 1947
`define FP16_TO_INDEX_3B4E 1948
`define FP16_TO_INDEX_3B52 1949
`define FP16_TO_INDEX_3B56 1950
`define FP16_TO_INDEX_3B5A 1951
`define FP16_TO_INDEX_3B5E 1952
`define FP16_TO_INDEX_3B62 1953
`define FP16_TO_INDEX_3B66 1954
`define FP16_TO_INDEX_3B6B 1955
`define FP16_TO_INDEX_3B6F 1956
`define FP16_TO_INDEX_3B73 1957
`define FP16_TO_INDEX_3B77 1958
`define FP16_TO_INDEX_3B7B 1959
`define FP16_TO_INDEX_3B7F 1960
`define FP16_TO_INDEX_3B83 1961
`define FP16_TO_INDEX_3B87 1962
`define FP16_TO_INDEX_3B8B 1963
`define FP16_TO_INDEX_3B90 1964
`define FP16_TO_INDEX_3B94 1965
`define FP16_TO_INDEX_3B98 1966
`define FP16_TO_INDEX_3B9C 1967
`define FP16_TO_INDEX_3BA0 1968
`define FP16_TO_INDEX_3BA4 1969
`define FP16_TO_INDEX_3BA8 1970
`define FP16_TO_INDEX_3BAC 1971
`define FP16_TO_INDEX_3BB0 1972
`define FP16_TO_INDEX_3BB5 1973
`define FP16_TO_INDEX_3BB9 1974
`define FP16_TO_INDEX_3BBD 1975
`define FP16_TO_INDEX_3BC1 1976
`define FP16_TO_INDEX_3BC5 1977
`define FP16_TO_INDEX_3BC9 1978
`define FP16_TO_INDEX_3BCD 1979
`define FP16_TO_INDEX_3BD1 1980
`define FP16_TO_INDEX_3BD5 1981
`define FP16_TO_INDEX_3BDA 1982
`define FP16_TO_INDEX_3BDE 1983
`define FP16_TO_INDEX_3BE2 1984
`define FP16_TO_INDEX_3BE6 1985
`define FP16_TO_INDEX_3BEA 1986
`define FP16_TO_INDEX_3BEE 1987
`define FP16_TO_INDEX_3BF2 1988
`define FP16_TO_INDEX_3BF6 1989
`define FP16_TO_INDEX_3BFB 1990
`define FP16_TO_INDEX_3BFF 1991
`define FP16_TO_INDEX_3C01 1992
`define FP16_TO_INDEX_3C03 1993
`define FP16_TO_INDEX_3C05 1994
`define FP16_TO_INDEX_3C08 1995
`define FP16_TO_INDEX_3C0A 1996
`define FP16_TO_INDEX_3C0C 1997
`define FP16_TO_INDEX_3C0E 1998
`define FP16_TO_INDEX_3C10 1999
`define FP16_TO_INDEX_3C12 2000
`define FP16_TO_INDEX_3C14 2001
`define FP16_TO_INDEX_3C16 2002
`define FP16_TO_INDEX_3C18 2003
`define FP16_TO_INDEX_3C1A 2004
`define FP16_TO_INDEX_3C1C 2005
`define FP16_TO_INDEX_3C1E 2006
`define FP16_TO_INDEX_3C20 2007
`define FP16_TO_INDEX_3C22 2008
`define FP16_TO_INDEX_3C24 2009
`define FP16_TO_INDEX_3C26 2010
`define FP16_TO_INDEX_3C28 2011
`define FP16_TO_INDEX_3C2B 2012
`define FP16_TO_INDEX_3C2D 2013
`define FP16_TO_INDEX_3C2F 2014
`define FP16_TO_INDEX_3C31 2015
`define FP16_TO_INDEX_3C33 2016
`define FP16_TO_INDEX_3C35 2017
`define FP16_TO_INDEX_3C37 2018
`define FP16_TO_INDEX_3C39 2019
`define FP16_TO_INDEX_3C3B 2020
`define FP16_TO_INDEX_3C3D 2021
`define FP16_TO_INDEX_3C3F 2022
`define FP16_TO_INDEX_3C41 2023
`define FP16_TO_INDEX_3C43 2024
`define FP16_TO_INDEX_3C45 2025
`define FP16_TO_INDEX_3C47 2026
`define FP16_TO_INDEX_3C49 2027
`define FP16_TO_INDEX_3C4B 2028
`define FP16_TO_INDEX_3C4D 2029
`define FP16_TO_INDEX_3C50 2030
`define FP16_TO_INDEX_3C52 2031
`define FP16_TO_INDEX_3C54 2032
`define FP16_TO_INDEX_3C56 2033
`define FP16_TO_INDEX_3C58 2034
`define FP16_TO_INDEX_3C5A 2035
`define FP16_TO_INDEX_3C5C 2036
`define FP16_TO_INDEX_3C5E 2037
`define FP16_TO_INDEX_3C60 2038
`define FP16_TO_INDEX_3C62 2039
`define FP16_TO_INDEX_3C64 2040
`define FP16_TO_INDEX_3C66 2041
`define FP16_TO_INDEX_3C68 2042
`define FP16_TO_INDEX_3C6A 2043
`define FP16_TO_INDEX_3C6C 2044
`define FP16_TO_INDEX_3C6E 2045
`define FP16_TO_INDEX_3C70 2046
`define FP16_TO_INDEX_3C73 2047
`define FP16_TO_INDEX_3C75 2048
`define FP16_TO_INDEX_3C77 2049
`define FP16_TO_INDEX_3C79 2050
`define FP16_TO_INDEX_3C7B 2051
`define FP16_TO_INDEX_3C7D 2052
`define FP16_TO_INDEX_3C7F 2053
`define FP16_TO_INDEX_3C81 2054
`define FP16_TO_INDEX_3C83 2055
`define FP16_TO_INDEX_3C85 2056
`define FP16_TO_INDEX_3C87 2057
`define FP16_TO_INDEX_3C89 2058
`define FP16_TO_INDEX_3C8B 2059
`define FP16_TO_INDEX_3C8D 2060
`define FP16_TO_INDEX_3C8F 2061
`define FP16_TO_INDEX_3C91 2062
`define FP16_TO_INDEX_3C93 2063
`define FP16_TO_INDEX_3C95 2064
`define FP16_TO_INDEX_3C98 2065
`define FP16_TO_INDEX_3C9A 2066
`define FP16_TO_INDEX_3C9C 2067
`define FP16_TO_INDEX_3C9E 2068
`define FP16_TO_INDEX_3CA0 2069
`define FP16_TO_INDEX_3CA2 2070
`define FP16_TO_INDEX_3CA4 2071
`define FP16_TO_INDEX_3CA6 2072
`define FP16_TO_INDEX_3CA8 2073
`define FP16_TO_INDEX_3CAA 2074
`define FP16_TO_INDEX_3CAC 2075
`define FP16_TO_INDEX_3CAE 2076
`define FP16_TO_INDEX_3CB0 2077
`define FP16_TO_INDEX_3CB2 2078
`define FP16_TO_INDEX_3CB4 2079
`define FP16_TO_INDEX_3CB6 2080
`define FP16_TO_INDEX_3CB8 2081
`define FP16_TO_INDEX_3CBA 2082
`define FP16_TO_INDEX_3CBD 2083
`define FP16_TO_INDEX_3CBF 2084
`define FP16_TO_INDEX_3CC1 2085
`define FP16_TO_INDEX_3CC3 2086
`define FP16_TO_INDEX_3CC5 2087
`define FP16_TO_INDEX_3CC7 2088
`define FP16_TO_INDEX_3CC9 2089
`define FP16_TO_INDEX_3CCB 2090
`define FP16_TO_INDEX_3CCD 2091
`define FP16_TO_INDEX_3CCF 2092
`define FP16_TO_INDEX_3CD1 2093
`define FP16_TO_INDEX_3CD3 2094
`define FP16_TO_INDEX_3CD5 2095
`define FP16_TO_INDEX_3CD7 2096
`define FP16_TO_INDEX_3CD9 2097
`define FP16_TO_INDEX_3CDB 2098
`define FP16_TO_INDEX_3CDD 2099
`define FP16_TO_INDEX_3CE0 2100
`define FP16_TO_INDEX_3CE2 2101
`define FP16_TO_INDEX_3CE4 2102
`define FP16_TO_INDEX_3CE6 2103
`define FP16_TO_INDEX_3CE8 2104
`define FP16_TO_INDEX_3CEA 2105
`define FP16_TO_INDEX_3CEC 2106
`define FP16_TO_INDEX_3CEE 2107
`define FP16_TO_INDEX_3CF0 2108
`define FP16_TO_INDEX_3CF2 2109
`define FP16_TO_INDEX_3CF4 2110
`define FP16_TO_INDEX_3CF6 2111
`define FP16_TO_INDEX_3CF8 2112
`define FP16_TO_INDEX_3CFA 2113
`define FP16_TO_INDEX_3CFC 2114
`define FP16_TO_INDEX_3CFE 2115
`define FP16_TO_INDEX_3D00 2116
`define FP16_TO_INDEX_3D02 2117
`define FP16_TO_INDEX_3D05 2118
`define FP16_TO_INDEX_3D07 2119
`define FP16_TO_INDEX_3D09 2120
`define FP16_TO_INDEX_3D0B 2121
`define FP16_TO_INDEX_3D0D 2122
`define FP16_TO_INDEX_3D0F 2123
`define FP16_TO_INDEX_3D11 2124
`define FP16_TO_INDEX_3D13 2125
`define FP16_TO_INDEX_3D15 2126
`define FP16_TO_INDEX_3D17 2127
`define FP16_TO_INDEX_3D19 2128
`define FP16_TO_INDEX_3D1B 2129
`define FP16_TO_INDEX_3D1D 2130
`define FP16_TO_INDEX_3D1F 2131
`define FP16_TO_INDEX_3D21 2132
`define FP16_TO_INDEX_3D23 2133
`define FP16_TO_INDEX_3D25 2134
`define FP16_TO_INDEX_3D28 2135
`define FP16_TO_INDEX_3D2A 2136
`define FP16_TO_INDEX_3D2C 2137
`define FP16_TO_INDEX_3D2E 2138
`define FP16_TO_INDEX_3D30 2139
`define FP16_TO_INDEX_3D32 2140
`define FP16_TO_INDEX_3D34 2141
`define FP16_TO_INDEX_3D36 2142
`define FP16_TO_INDEX_3D38 2143
`define FP16_TO_INDEX_3D3A 2144
`define FP16_TO_INDEX_3D3C 2145
`define FP16_TO_INDEX_3D3E 2146
`define FP16_TO_INDEX_3D40 2147
`define FP16_TO_INDEX_3D42 2148
`define FP16_TO_INDEX_3D44 2149
`define FP16_TO_INDEX_3D46 2150
`define FP16_TO_INDEX_3D48 2151
`define FP16_TO_INDEX_3D4A 2152
`define FP16_TO_INDEX_3D4D 2153
`define FP16_TO_INDEX_3D4F 2154
`define FP16_TO_INDEX_3D51 2155
`define FP16_TO_INDEX_3D53 2156
`define FP16_TO_INDEX_3D55 2157
`define FP16_TO_INDEX_3D57 2158
`define FP16_TO_INDEX_3D59 2159
`define FP16_TO_INDEX_3D5B 2160
`define FP16_TO_INDEX_3D5D 2161
`define FP16_TO_INDEX_3D5F 2162
`define FP16_TO_INDEX_3D61 2163
`define FP16_TO_INDEX_3D63 2164
`define FP16_TO_INDEX_3D65 2165
`define FP16_TO_INDEX_3D67 2166
`define FP16_TO_INDEX_3D69 2167
`define FP16_TO_INDEX_3D6B 2168
`define FP16_TO_INDEX_3D6D 2169
`define FP16_TO_INDEX_3D70 2170
`define FP16_TO_INDEX_3D72 2171
`define FP16_TO_INDEX_3D74 2172
`define FP16_TO_INDEX_3D76 2173
`define FP16_TO_INDEX_3D78 2174
`define FP16_TO_INDEX_3D7A 2175
`define FP16_TO_INDEX_3D7C 2176
`define FP16_TO_INDEX_3D7E 2177
`define FP16_TO_INDEX_3D80 2178
`define FP16_TO_INDEX_3D82 2179
`define FP16_TO_INDEX_3D84 2180
`define FP16_TO_INDEX_3D86 2181
`define FP16_TO_INDEX_3D88 2182
`define FP16_TO_INDEX_3D8A 2183
`define FP16_TO_INDEX_3D8C 2184
`define FP16_TO_INDEX_3D8E 2185
`define FP16_TO_INDEX_3D90 2186
`define FP16_TO_INDEX_3D92 2187
`define FP16_TO_INDEX_3D95 2188
`define FP16_TO_INDEX_3D97 2189
`define FP16_TO_INDEX_3D99 2190
`define FP16_TO_INDEX_3D9B 2191
`define FP16_TO_INDEX_3D9D 2192
`define FP16_TO_INDEX_3D9F 2193
`define FP16_TO_INDEX_3DA1 2194
`define FP16_TO_INDEX_3DA3 2195
`define FP16_TO_INDEX_3DA5 2196
`define FP16_TO_INDEX_3DA7 2197
`define FP16_TO_INDEX_3DA9 2198
`define FP16_TO_INDEX_3DAB 2199
`define FP16_TO_INDEX_3DAD 2200
`define FP16_TO_INDEX_3DAF 2201
`define FP16_TO_INDEX_3DB1 2202
`define FP16_TO_INDEX_3DB3 2203
`define FP16_TO_INDEX_3DB5 2204
`define FP16_TO_INDEX_3DB7 2205
`define FP16_TO_INDEX_3DBA 2206
`define FP16_TO_INDEX_3DBC 2207
`define FP16_TO_INDEX_3DBE 2208
`define FP16_TO_INDEX_3DC0 2209
`define FP16_TO_INDEX_3DC2 2210
`define FP16_TO_INDEX_3DC4 2211
`define FP16_TO_INDEX_3DC6 2212
`define FP16_TO_INDEX_3DC8 2213
`define FP16_TO_INDEX_3DCA 2214
`define FP16_TO_INDEX_3DCC 2215
`define FP16_TO_INDEX_3DCE 2216
`define FP16_TO_INDEX_3DD0 2217
`define FP16_TO_INDEX_3DD2 2218
`define FP16_TO_INDEX_3DD4 2219
`define FP16_TO_INDEX_3DD6 2220
`define FP16_TO_INDEX_3DD8 2221
`define FP16_TO_INDEX_3DDA 2222
`define FP16_TO_INDEX_3DDD 2223
`define FP16_TO_INDEX_3DDF 2224
`define FP16_TO_INDEX_3DE1 2225
`define FP16_TO_INDEX_3DE3 2226
`define FP16_TO_INDEX_3DE5 2227
`define FP16_TO_INDEX_3DE7 2228
`define FP16_TO_INDEX_3DE9 2229
`define FP16_TO_INDEX_3DEB 2230
`define FP16_TO_INDEX_3DED 2231
`define FP16_TO_INDEX_3DEF 2232
`define FP16_TO_INDEX_3DF1 2233
`define FP16_TO_INDEX_3DF3 2234
`define FP16_TO_INDEX_3DF5 2235
`define FP16_TO_INDEX_3DF7 2236
`define FP16_TO_INDEX_3DF9 2237
`define FP16_TO_INDEX_3DFB 2238
`define FP16_TO_INDEX_3DFD 2239
`define FP16_TO_INDEX_3DFF 2240
`define FP16_TO_INDEX_3E02 2241
`define FP16_TO_INDEX_3E04 2242
`define FP16_TO_INDEX_3E06 2243
`define FP16_TO_INDEX_3E08 2244
`define FP16_TO_INDEX_3E0A 2245
`define FP16_TO_INDEX_3E0C 2246
`define FP16_TO_INDEX_3E0E 2247
`define FP16_TO_INDEX_3E10 2248
`define FP16_TO_INDEX_3E12 2249
`define FP16_TO_INDEX_3E14 2250
`define FP16_TO_INDEX_3E16 2251
`define FP16_TO_INDEX_3E18 2252
`define FP16_TO_INDEX_3E1A 2253
`define FP16_TO_INDEX_3E1C 2254
`define FP16_TO_INDEX_3E1E 2255
`define FP16_TO_INDEX_3E20 2256
`define FP16_TO_INDEX_3E22 2257
`define FP16_TO_INDEX_3E25 2258
`define FP16_TO_INDEX_3E27 2259
`define FP16_TO_INDEX_3E29 2260
`define FP16_TO_INDEX_3E2B 2261
`define FP16_TO_INDEX_3E2D 2262
`define FP16_TO_INDEX_3E2F 2263
`define FP16_TO_INDEX_3E31 2264
`define FP16_TO_INDEX_3E33 2265
`define FP16_TO_INDEX_3E35 2266
`define FP16_TO_INDEX_3E37 2267
`define FP16_TO_INDEX_3E39 2268
`define FP16_TO_INDEX_3E3B 2269
`define FP16_TO_INDEX_3E3D 2270
`define FP16_TO_INDEX_3E3F 2271
`define FP16_TO_INDEX_3E41 2272
`define FP16_TO_INDEX_3E43 2273
`define FP16_TO_INDEX_3E45 2274
`define FP16_TO_INDEX_3E47 2275
`define FP16_TO_INDEX_3E4A 2276
`define FP16_TO_INDEX_3E4C 2277
`define FP16_TO_INDEX_3E4E 2278
`define FP16_TO_INDEX_3E50 2279
`define FP16_TO_INDEX_3E52 2280
`define FP16_TO_INDEX_3E54 2281
`define FP16_TO_INDEX_3E56 2282
`define FP16_TO_INDEX_3E58 2283
`define FP16_TO_INDEX_3E5A 2284
`define FP16_TO_INDEX_3E5C 2285
`define FP16_TO_INDEX_3E5E 2286
`define FP16_TO_INDEX_3E60 2287
`define FP16_TO_INDEX_3E62 2288
`define FP16_TO_INDEX_3E64 2289
`define FP16_TO_INDEX_3E66 2290
`define FP16_TO_INDEX_3E68 2291
`define FP16_TO_INDEX_3E6A 2292
`define FP16_TO_INDEX_3E6D 2293
`define FP16_TO_INDEX_3E6F 2294
`define FP16_TO_INDEX_3E71 2295
`define FP16_TO_INDEX_3E73 2296
`define FP16_TO_INDEX_3E75 2297
`define FP16_TO_INDEX_3E77 2298
`define FP16_TO_INDEX_3E79 2299
`define FP16_TO_INDEX_3E7B 2300
`define FP16_TO_INDEX_3E7D 2301
`define FP16_TO_INDEX_3E7F 2302
`define FP16_TO_INDEX_3E81 2303
`define FP16_TO_INDEX_3E83 2304
`define FP16_TO_INDEX_3E85 2305
`define FP16_TO_INDEX_3E87 2306
`define FP16_TO_INDEX_3E89 2307
`define FP16_TO_INDEX_3E8B 2308
`define FP16_TO_INDEX_3E8D 2309
`define FP16_TO_INDEX_3E8F 2310
`define FP16_TO_INDEX_3E92 2311
`define FP16_TO_INDEX_3E94 2312
`define FP16_TO_INDEX_3E96 2313
`define FP16_TO_INDEX_3E98 2314
`define FP16_TO_INDEX_3E9A 2315
`define FP16_TO_INDEX_3E9C 2316
`define FP16_TO_INDEX_3E9E 2317
`define FP16_TO_INDEX_3EA0 2318
`define FP16_TO_INDEX_3EA2 2319
`define FP16_TO_INDEX_3EA4 2320
`define FP16_TO_INDEX_3EA6 2321
`define FP16_TO_INDEX_3EA8 2322
`define FP16_TO_INDEX_3EAA 2323
`define FP16_TO_INDEX_3EAC 2324
`define FP16_TO_INDEX_3EAE 2325
`define FP16_TO_INDEX_3EB0 2326
`define FP16_TO_INDEX_3EB2 2327
`define FP16_TO_INDEX_3EB4 2328
`define FP16_TO_INDEX_3EB7 2329
`define FP16_TO_INDEX_3EB9 2330
`define FP16_TO_INDEX_3EBB 2331
`define FP16_TO_INDEX_3EBD 2332
`define FP16_TO_INDEX_3EBF 2333
`define FP16_TO_INDEX_3EC1 2334
`define FP16_TO_INDEX_3EC3 2335
`define FP16_TO_INDEX_3EC5 2336
`define FP16_TO_INDEX_3EC7 2337
`define FP16_TO_INDEX_3EC9 2338
`define FP16_TO_INDEX_3ECB 2339
`define FP16_TO_INDEX_3ECD 2340
`define FP16_TO_INDEX_3ECF 2341
`define FP16_TO_INDEX_3ED1 2342
`define FP16_TO_INDEX_3ED3 2343
`define FP16_TO_INDEX_3ED5 2344
`define FP16_TO_INDEX_3ED7 2345
`define FP16_TO_INDEX_3EDA 2346
`define FP16_TO_INDEX_3EDC 2347
`define FP16_TO_INDEX_3EDE 2348
`define FP16_TO_INDEX_3EE0 2349
`define FP16_TO_INDEX_3EE2 2350
`define FP16_TO_INDEX_3EE4 2351
`define FP16_TO_INDEX_3EE6 2352
`define FP16_TO_INDEX_3EE8 2353
`define FP16_TO_INDEX_3EEA 2354
`define FP16_TO_INDEX_3EEC 2355
`define FP16_TO_INDEX_3EEE 2356
`define FP16_TO_INDEX_3EF0 2357
`define FP16_TO_INDEX_3EF2 2358
`define FP16_TO_INDEX_3EF4 2359
`define FP16_TO_INDEX_3EF6 2360
`define FP16_TO_INDEX_3EF8 2361
`define FP16_TO_INDEX_3EFA 2362
`define FP16_TO_INDEX_3EFC 2363
`define FP16_TO_INDEX_3EFF 2364
`define FP16_TO_INDEX_3F01 2365
`define FP16_TO_INDEX_3F03 2366
`define FP16_TO_INDEX_3F05 2367
`define FP16_TO_INDEX_3F07 2368
`define FP16_TO_INDEX_3F09 2369
`define FP16_TO_INDEX_3F0B 2370
`define FP16_TO_INDEX_3F0D 2371
`define FP16_TO_INDEX_3F0F 2372
`define FP16_TO_INDEX_3F11 2373
`define FP16_TO_INDEX_3F13 2374
`define FP16_TO_INDEX_3F15 2375
`define FP16_TO_INDEX_3F17 2376
`define FP16_TO_INDEX_3F19 2377
`define FP16_TO_INDEX_3F1B 2378
`define FP16_TO_INDEX_3F1D 2379
`define FP16_TO_INDEX_3F1F 2380
`define FP16_TO_INDEX_3F22 2381
`define FP16_TO_INDEX_3F24 2382
`define FP16_TO_INDEX_3F26 2383
`define FP16_TO_INDEX_3F28 2384
`define FP16_TO_INDEX_3F2A 2385
`define FP16_TO_INDEX_3F2C 2386
`define FP16_TO_INDEX_3F2E 2387
`define FP16_TO_INDEX_3F30 2388
`define FP16_TO_INDEX_3F32 2389
`define FP16_TO_INDEX_3F34 2390
`define FP16_TO_INDEX_3F36 2391
`define FP16_TO_INDEX_3F38 2392
`define FP16_TO_INDEX_3F3A 2393
`define FP16_TO_INDEX_3F3C 2394
`define FP16_TO_INDEX_3F3E 2395
`define FP16_TO_INDEX_3F40 2396
`define FP16_TO_INDEX_3F42 2397
`define FP16_TO_INDEX_3F44 2398
`define FP16_TO_INDEX_3F47 2399
`define FP16_TO_INDEX_3F49 2400
`define FP16_TO_INDEX_3F4B 2401
`define FP16_TO_INDEX_3F4D 2402
`define FP16_TO_INDEX_3F4F 2403
`define FP16_TO_INDEX_3F51 2404
`define FP16_TO_INDEX_3F53 2405
`define FP16_TO_INDEX_3F55 2406
`define FP16_TO_INDEX_3F57 2407
`define FP16_TO_INDEX_3F59 2408
`define FP16_TO_INDEX_3F5B 2409
`define FP16_TO_INDEX_3F5D 2410
`define FP16_TO_INDEX_3F5F 2411
`define FP16_TO_INDEX_3F61 2412
`define FP16_TO_INDEX_3F63 2413
`define FP16_TO_INDEX_3F65 2414
`define FP16_TO_INDEX_3F67 2415
`define FP16_TO_INDEX_3F6A 2416
`define FP16_TO_INDEX_3F6C 2417
`define FP16_TO_INDEX_3F6E 2418
`define FP16_TO_INDEX_3F70 2419
`define FP16_TO_INDEX_3F72 2420
`define FP16_TO_INDEX_3F74 2421
`define FP16_TO_INDEX_3F76 2422
`define FP16_TO_INDEX_3F78 2423
`define FP16_TO_INDEX_3F7A 2424
`define FP16_TO_INDEX_3F7C 2425
`define FP16_TO_INDEX_3F7E 2426
`define FP16_TO_INDEX_3F80 2427
`define FP16_TO_INDEX_3F82 2428
`define FP16_TO_INDEX_3F84 2429
`define FP16_TO_INDEX_3F86 2430
`define FP16_TO_INDEX_3F88 2431
`define FP16_TO_INDEX_3F8A 2432
`define FP16_TO_INDEX_3F8C 2433
`define FP16_TO_INDEX_3F8F 2434
`define FP16_TO_INDEX_3F91 2435
`define FP16_TO_INDEX_3F93 2436
`define FP16_TO_INDEX_3F95 2437
`define FP16_TO_INDEX_3F97 2438
`define FP16_TO_INDEX_3F99 2439
`define FP16_TO_INDEX_3F9B 2440
`define FP16_TO_INDEX_3F9D 2441
`define FP16_TO_INDEX_3F9F 2442
`define FP16_TO_INDEX_3FA1 2443
`define FP16_TO_INDEX_3FA3 2444
`define FP16_TO_INDEX_3FA5 2445
`define FP16_TO_INDEX_3FA7 2446
`define FP16_TO_INDEX_3FA9 2447
`define FP16_TO_INDEX_3FAB 2448
`define FP16_TO_INDEX_3FAD 2449
`define FP16_TO_INDEX_3FAF 2450
`define FP16_TO_INDEX_3FB1 2451
`define FP16_TO_INDEX_3FB4 2452
`define FP16_TO_INDEX_3FB6 2453
`define FP16_TO_INDEX_3FB8 2454
`define FP16_TO_INDEX_3FBA 2455
`define FP16_TO_INDEX_3FBC 2456
`define FP16_TO_INDEX_3FBE 2457
`define FP16_TO_INDEX_3FC0 2458
`define FP16_TO_INDEX_3FC2 2459
`define FP16_TO_INDEX_3FC4 2460
`define FP16_TO_INDEX_3FC6 2461
`define FP16_TO_INDEX_3FC8 2462
`define FP16_TO_INDEX_3FCA 2463
`define FP16_TO_INDEX_3FCC 2464
`define FP16_TO_INDEX_3FCE 2465
`define FP16_TO_INDEX_3FD0 2466
`define FP16_TO_INDEX_3FD2 2467
`define FP16_TO_INDEX_3FD4 2468
`define FP16_TO_INDEX_3FD7 2469
`define FP16_TO_INDEX_3FD9 2470
`define FP16_TO_INDEX_3FDB 2471
`define FP16_TO_INDEX_3FDD 2472
`define FP16_TO_INDEX_3FDF 2473
`define FP16_TO_INDEX_3FE1 2474
`define FP16_TO_INDEX_3FE3 2475
`define FP16_TO_INDEX_3FE5 2476
`define FP16_TO_INDEX_3FE7 2477
`define FP16_TO_INDEX_3FE9 2478
`define FP16_TO_INDEX_3FEB 2479
`define FP16_TO_INDEX_3FED 2480
`define FP16_TO_INDEX_3FEF 2481
`define FP16_TO_INDEX_3FF1 2482
`define FP16_TO_INDEX_3FF3 2483
`define FP16_TO_INDEX_3FF5 2484
`define FP16_TO_INDEX_3FF7 2485
`define FP16_TO_INDEX_3FF9 2486
`define FP16_TO_INDEX_3FFC 2487
`define FP16_TO_INDEX_3FFE 2488
`define FP16_TO_INDEX_4000 2489
`define FP16_TO_INDEX_4001 2490
`define FP16_TO_INDEX_4002 2491
`define FP16_TO_INDEX_4003 2492
`define FP16_TO_INDEX_4004 2493
`define FP16_TO_INDEX_4005 2494
`define FP16_TO_INDEX_4006 2495
`define FP16_TO_INDEX_4007 2496
`define FP16_TO_INDEX_4008 2497
`define FP16_TO_INDEX_4009 2498
`define FP16_TO_INDEX_400A 2499
`define FP16_TO_INDEX_400B 2500
`define FP16_TO_INDEX_400C 2501
`define FP16_TO_INDEX_400D 2502
`define FP16_TO_INDEX_400E 2503
`define FP16_TO_INDEX_400F 2504
`define FP16_TO_INDEX_4010 2505
`define FP16_TO_INDEX_4011 2506
`define FP16_TO_INDEX_4012 2507
`define FP16_TO_INDEX_4013 2508
`define FP16_TO_INDEX_4014 2509
`define FP16_TO_INDEX_4015 2510
`define FP16_TO_INDEX_4016 2511
`define FP16_TO_INDEX_4017 2512
`define FP16_TO_INDEX_4019 2513
`define FP16_TO_INDEX_401A 2514
`define FP16_TO_INDEX_401B 2515
`define FP16_TO_INDEX_401C 2516
`define FP16_TO_INDEX_401D 2517
`define FP16_TO_INDEX_401E 2518
`define FP16_TO_INDEX_401F 2519
`define FP16_TO_INDEX_4020 2520
`define FP16_TO_INDEX_4021 2521
`define FP16_TO_INDEX_4022 2522
`define FP16_TO_INDEX_4023 2523
`define FP16_TO_INDEX_4024 2524
`define FP16_TO_INDEX_4025 2525
`define FP16_TO_INDEX_4026 2526
`define FP16_TO_INDEX_4027 2527
`define FP16_TO_INDEX_4028 2528
`define FP16_TO_INDEX_4029 2529
`define FP16_TO_INDEX_402A 2530
`define FP16_TO_INDEX_402B 2531
`define FP16_TO_INDEX_402C 2532
`define FP16_TO_INDEX_402D 2533
`define FP16_TO_INDEX_402E 2534
`define FP16_TO_INDEX_402F 2535
`define FP16_TO_INDEX_4030 2536
`define FP16_TO_INDEX_4031 2537
`define FP16_TO_INDEX_4032 2538
`define FP16_TO_INDEX_4033 2539
`define FP16_TO_INDEX_4034 2540
`define FP16_TO_INDEX_4035 2541
`define FP16_TO_INDEX_4036 2542
`define FP16_TO_INDEX_4037 2543
`define FP16_TO_INDEX_4038 2544
`define FP16_TO_INDEX_4039 2545
`define FP16_TO_INDEX_403A 2546
`define FP16_TO_INDEX_403B 2547
`define FP16_TO_INDEX_403D 2548
`define FP16_TO_INDEX_403E 2549
`define FP16_TO_INDEX_403F 2550
`define FP16_TO_INDEX_4040 2551
`define FP16_TO_INDEX_4041 2552
`define FP16_TO_INDEX_4042 2553
`define FP16_TO_INDEX_4043 2554
`define FP16_TO_INDEX_4044 2555
`define FP16_TO_INDEX_4045 2556
`define FP16_TO_INDEX_4046 2557
`define FP16_TO_INDEX_4047 2558
`define FP16_TO_INDEX_4048 2559
`define FP16_TO_INDEX_4049 2560
`define FP16_TO_INDEX_404A 2561
`define FP16_TO_INDEX_404B 2562
`define FP16_TO_INDEX_404C 2563
`define FP16_TO_INDEX_404D 2564
`define FP16_TO_INDEX_404E 2565
`define FP16_TO_INDEX_404F 2566
`define FP16_TO_INDEX_4050 2567
`define FP16_TO_INDEX_4051 2568
`define FP16_TO_INDEX_4052 2569
`define FP16_TO_INDEX_4053 2570
`define FP16_TO_INDEX_4054 2571
`define FP16_TO_INDEX_4055 2572
`define FP16_TO_INDEX_4056 2573
`define FP16_TO_INDEX_4057 2574
`define FP16_TO_INDEX_4058 2575
`define FP16_TO_INDEX_4059 2576
`define FP16_TO_INDEX_405A 2577
`define FP16_TO_INDEX_405B 2578
`define FP16_TO_INDEX_405C 2579
`define FP16_TO_INDEX_405D 2580
`define FP16_TO_INDEX_405E 2581
`define FP16_TO_INDEX_405F 2582
`define FP16_TO_INDEX_4061 2583
`define FP16_TO_INDEX_4062 2584
`define FP16_TO_INDEX_4063 2585
`define FP16_TO_INDEX_4064 2586
`define FP16_TO_INDEX_4065 2587
`define FP16_TO_INDEX_4066 2588
`define FP16_TO_INDEX_4067 2589
`define FP16_TO_INDEX_4068 2590
`define FP16_TO_INDEX_4069 2591
`define FP16_TO_INDEX_406A 2592
`define FP16_TO_INDEX_406B 2593
`define FP16_TO_INDEX_406C 2594
`define FP16_TO_INDEX_406D 2595
`define FP16_TO_INDEX_406E 2596
`define FP16_TO_INDEX_406F 2597
`define FP16_TO_INDEX_4070 2598
`define FP16_TO_INDEX_4071 2599
`define FP16_TO_INDEX_4072 2600
`define FP16_TO_INDEX_4073 2601
`define FP16_TO_INDEX_4074 2602
`define FP16_TO_INDEX_4075 2603
`define FP16_TO_INDEX_4076 2604
`define FP16_TO_INDEX_4077 2605
`define FP16_TO_INDEX_4078 2606
`define FP16_TO_INDEX_4079 2607
`define FP16_TO_INDEX_407A 2608
`define FP16_TO_INDEX_407B 2609
`define FP16_TO_INDEX_407C 2610
`define FP16_TO_INDEX_407D 2611
`define FP16_TO_INDEX_407E 2612
`define FP16_TO_INDEX_407F 2613
`define FP16_TO_INDEX_4080 2614
`define FP16_TO_INDEX_4081 2615
`define FP16_TO_INDEX_4082 2616
`define FP16_TO_INDEX_4083 2617
`define FP16_TO_INDEX_4084 2618
`define FP16_TO_INDEX_4086 2619
`define FP16_TO_INDEX_4087 2620
`define FP16_TO_INDEX_4088 2621
`define FP16_TO_INDEX_4089 2622
`define FP16_TO_INDEX_408A 2623
`define FP16_TO_INDEX_408B 2624
`define FP16_TO_INDEX_408C 2625
`define FP16_TO_INDEX_408D 2626
`define FP16_TO_INDEX_408E 2627
`define FP16_TO_INDEX_408F 2628
`define FP16_TO_INDEX_4090 2629
`define FP16_TO_INDEX_4091 2630
`define FP16_TO_INDEX_4092 2631
`define FP16_TO_INDEX_4093 2632
`define FP16_TO_INDEX_4094 2633
`define FP16_TO_INDEX_4095 2634
`define FP16_TO_INDEX_4096 2635
`define FP16_TO_INDEX_4097 2636
`define FP16_TO_INDEX_4098 2637
`define FP16_TO_INDEX_4099 2638
`define FP16_TO_INDEX_409A 2639
`define FP16_TO_INDEX_409B 2640
`define FP16_TO_INDEX_409C 2641
`define FP16_TO_INDEX_409D 2642
`define FP16_TO_INDEX_409E 2643
`define FP16_TO_INDEX_409F 2644
`define FP16_TO_INDEX_40A0 2645
`define FP16_TO_INDEX_40A1 2646
`define FP16_TO_INDEX_40A2 2647
`define FP16_TO_INDEX_40A3 2648
`define FP16_TO_INDEX_40A4 2649
`define FP16_TO_INDEX_40A5 2650
`define FP16_TO_INDEX_40A6 2651
`define FP16_TO_INDEX_40A7 2652
`define FP16_TO_INDEX_40A8 2653
`define FP16_TO_INDEX_40AA 2654
`define FP16_TO_INDEX_40AB 2655
`define FP16_TO_INDEX_40AC 2656
`define FP16_TO_INDEX_40AD 2657
`define FP16_TO_INDEX_40AE 2658
`define FP16_TO_INDEX_40AF 2659
`define FP16_TO_INDEX_40B0 2660
`define FP16_TO_INDEX_40B1 2661
`define FP16_TO_INDEX_40B2 2662
`define FP16_TO_INDEX_40B3 2663
`define FP16_TO_INDEX_40B4 2664
`define FP16_TO_INDEX_40B5 2665
`define FP16_TO_INDEX_40B6 2666
`define FP16_TO_INDEX_40B7 2667
`define FP16_TO_INDEX_40B8 2668
`define FP16_TO_INDEX_40B9 2669
`define FP16_TO_INDEX_40BA 2670
`define FP16_TO_INDEX_40BB 2671
`define FP16_TO_INDEX_40BC 2672
`define FP16_TO_INDEX_40BD 2673
`define FP16_TO_INDEX_40BE 2674
`define FP16_TO_INDEX_40BF 2675
`define FP16_TO_INDEX_40C0 2676
`define FP16_TO_INDEX_40C1 2677
`define FP16_TO_INDEX_40C2 2678
`define FP16_TO_INDEX_40C3 2679
`define FP16_TO_INDEX_40C4 2680
`define FP16_TO_INDEX_40C5 2681
`define FP16_TO_INDEX_40C6 2682
`define FP16_TO_INDEX_40C7 2683
`define FP16_TO_INDEX_40C8 2684
`define FP16_TO_INDEX_40C9 2685
`define FP16_TO_INDEX_40CA 2686
`define FP16_TO_INDEX_40CB 2687
`define FP16_TO_INDEX_40CC 2688
`define FP16_TO_INDEX_40CE 2689
`define FP16_TO_INDEX_40CF 2690
`define FP16_TO_INDEX_40D0 2691
`define FP16_TO_INDEX_40D1 2692
`define FP16_TO_INDEX_40D2 2693
`define FP16_TO_INDEX_40D3 2694
`define FP16_TO_INDEX_40D4 2695
`define FP16_TO_INDEX_40D5 2696
`define FP16_TO_INDEX_40D6 2697
`define FP16_TO_INDEX_40D7 2698
`define FP16_TO_INDEX_40D8 2699
`define FP16_TO_INDEX_40D9 2700
`define FP16_TO_INDEX_40DA 2701
`define FP16_TO_INDEX_40DB 2702
`define FP16_TO_INDEX_40DC 2703
`define FP16_TO_INDEX_40DD 2704
`define FP16_TO_INDEX_40DE 2705
`define FP16_TO_INDEX_40DF 2706
`define FP16_TO_INDEX_40E0 2707
`define FP16_TO_INDEX_40E1 2708
`define FP16_TO_INDEX_40E2 2709
`define FP16_TO_INDEX_40E3 2710
`define FP16_TO_INDEX_40E4 2711
`define FP16_TO_INDEX_40E5 2712
`define FP16_TO_INDEX_40E6 2713
`define FP16_TO_INDEX_40E7 2714
`define FP16_TO_INDEX_40E8 2715
`define FP16_TO_INDEX_40E9 2716
`define FP16_TO_INDEX_40EA 2717
`define FP16_TO_INDEX_40EB 2718
`define FP16_TO_INDEX_40EC 2719
`define FP16_TO_INDEX_40ED 2720
`define FP16_TO_INDEX_40EE 2721
`define FP16_TO_INDEX_40EF 2722
`define FP16_TO_INDEX_40F0 2723
`define FP16_TO_INDEX_40F2 2724
`define FP16_TO_INDEX_40F3 2725
`define FP16_TO_INDEX_40F4 2726
`define FP16_TO_INDEX_40F5 2727
`define FP16_TO_INDEX_40F6 2728
`define FP16_TO_INDEX_40F7 2729
`define FP16_TO_INDEX_40F8 2730
`define FP16_TO_INDEX_40F9 2731
`define FP16_TO_INDEX_40FA 2732
`define FP16_TO_INDEX_40FB 2733
`define FP16_TO_INDEX_40FC 2734
`define FP16_TO_INDEX_40FD 2735
`define FP16_TO_INDEX_40FE 2736
`define FP16_TO_INDEX_40FF 2737
`define FP16_TO_INDEX_4100 2738
`define FP16_TO_INDEX_4101 2739
`define FP16_TO_INDEX_4102 2740
`define FP16_TO_INDEX_4103 2741
`define FP16_TO_INDEX_4104 2742
`define FP16_TO_INDEX_4105 2743
`define FP16_TO_INDEX_4106 2744
`define FP16_TO_INDEX_4107 2745
`define FP16_TO_INDEX_4108 2746
`define FP16_TO_INDEX_4109 2747
`define FP16_TO_INDEX_410A 2748
`define FP16_TO_INDEX_410B 2749
`define FP16_TO_INDEX_410C 2750
`define FP16_TO_INDEX_410D 2751
`define FP16_TO_INDEX_410E 2752
`define FP16_TO_INDEX_410F 2753
`define FP16_TO_INDEX_4110 2754
`define FP16_TO_INDEX_4111 2755
`define FP16_TO_INDEX_4112 2756
`define FP16_TO_INDEX_4113 2757
`define FP16_TO_INDEX_4114 2758
`define FP16_TO_INDEX_4116 2759
`define FP16_TO_INDEX_4117 2760
`define FP16_TO_INDEX_4118 2761
`define FP16_TO_INDEX_4119 2762
`define FP16_TO_INDEX_411A 2763
`define FP16_TO_INDEX_411B 2764
`define FP16_TO_INDEX_411C 2765
`define FP16_TO_INDEX_411D 2766
`define FP16_TO_INDEX_411E 2767
`define FP16_TO_INDEX_411F 2768
`define FP16_TO_INDEX_4120 2769
`define FP16_TO_INDEX_4121 2770
`define FP16_TO_INDEX_4122 2771
`define FP16_TO_INDEX_4123 2772
`define FP16_TO_INDEX_4124 2773
`define FP16_TO_INDEX_4125 2774
`define FP16_TO_INDEX_4126 2775
`define FP16_TO_INDEX_4127 2776
`define FP16_TO_INDEX_4128 2777
`define FP16_TO_INDEX_4129 2778
`define FP16_TO_INDEX_412A 2779
`define FP16_TO_INDEX_412B 2780
`define FP16_TO_INDEX_412C 2781
`define FP16_TO_INDEX_412D 2782
`define FP16_TO_INDEX_412E 2783
`define FP16_TO_INDEX_412F 2784
`define FP16_TO_INDEX_4130 2785
`define FP16_TO_INDEX_4131 2786
`define FP16_TO_INDEX_4132 2787
`define FP16_TO_INDEX_4133 2788
`define FP16_TO_INDEX_4134 2789
`define FP16_TO_INDEX_4135 2790
`define FP16_TO_INDEX_4136 2791
`define FP16_TO_INDEX_4137 2792
`define FP16_TO_INDEX_4138 2793
`define FP16_TO_INDEX_413A 2794
`define FP16_TO_INDEX_413B 2795
`define FP16_TO_INDEX_413C 2796
`define FP16_TO_INDEX_413D 2797
`define FP16_TO_INDEX_413E 2798
`define FP16_TO_INDEX_413F 2799
`define FP16_TO_INDEX_4140 2800
`define FP16_TO_INDEX_4141 2801
`define FP16_TO_INDEX_4142 2802
`define FP16_TO_INDEX_4143 2803
`define FP16_TO_INDEX_4144 2804
`define FP16_TO_INDEX_4145 2805
`define FP16_TO_INDEX_4146 2806
`define FP16_TO_INDEX_4147 2807
`define FP16_TO_INDEX_4148 2808
`define FP16_TO_INDEX_4149 2809
`define FP16_TO_INDEX_414A 2810
`define FP16_TO_INDEX_414B 2811
`define FP16_TO_INDEX_414C 2812
`define FP16_TO_INDEX_414D 2813
`define FP16_TO_INDEX_414E 2814
`define FP16_TO_INDEX_414F 2815
`define FP16_TO_INDEX_4150 2816
`define FP16_TO_INDEX_4151 2817
`define FP16_TO_INDEX_4152 2818
`define FP16_TO_INDEX_4153 2819
`define FP16_TO_INDEX_4154 2820
`define FP16_TO_INDEX_4155 2821
`define FP16_TO_INDEX_4156 2822
`define FP16_TO_INDEX_4157 2823
`define FP16_TO_INDEX_4158 2824
`define FP16_TO_INDEX_4159 2825
`define FP16_TO_INDEX_415A 2826
`define FP16_TO_INDEX_415B 2827
`define FP16_TO_INDEX_415C 2828
`define FP16_TO_INDEX_415E 2829
`define FP16_TO_INDEX_415F 2830
`define FP16_TO_INDEX_4160 2831
`define FP16_TO_INDEX_4161 2832
`define FP16_TO_INDEX_4162 2833
`define FP16_TO_INDEX_4163 2834
`define FP16_TO_INDEX_4164 2835
`define FP16_TO_INDEX_4165 2836
`define FP16_TO_INDEX_4166 2837
`define FP16_TO_INDEX_4167 2838
`define FP16_TO_INDEX_4168 2839
`define FP16_TO_INDEX_4169 2840
`define FP16_TO_INDEX_416A 2841
`define FP16_TO_INDEX_416B 2842
`define FP16_TO_INDEX_416C 2843
`define FP16_TO_INDEX_416D 2844
`define FP16_TO_INDEX_416E 2845
`define FP16_TO_INDEX_416F 2846
`define FP16_TO_INDEX_4170 2847
`define FP16_TO_INDEX_4171 2848
`define FP16_TO_INDEX_4172 2849
`define FP16_TO_INDEX_4173 2850
`define FP16_TO_INDEX_4174 2851
`define FP16_TO_INDEX_4175 2852
`define FP16_TO_INDEX_4176 2853
`define FP16_TO_INDEX_4177 2854
`define FP16_TO_INDEX_4178 2855
`define FP16_TO_INDEX_4179 2856
`define FP16_TO_INDEX_417A 2857
`define FP16_TO_INDEX_417B 2858
`define FP16_TO_INDEX_417C 2859
`define FP16_TO_INDEX_417D 2860
`define FP16_TO_INDEX_417E 2861
`define FP16_TO_INDEX_417F 2862
`define FP16_TO_INDEX_4180 2863
`define FP16_TO_INDEX_4181 2864
`define FP16_TO_INDEX_4183 2865
`define FP16_TO_INDEX_4184 2866
`define FP16_TO_INDEX_4185 2867
`define FP16_TO_INDEX_4186 2868
`define FP16_TO_INDEX_4187 2869
`define FP16_TO_INDEX_4188 2870
`define FP16_TO_INDEX_4189 2871
`define FP16_TO_INDEX_418A 2872
`define FP16_TO_INDEX_418B 2873
`define FP16_TO_INDEX_418C 2874
`define FP16_TO_INDEX_418D 2875
`define FP16_TO_INDEX_418E 2876
`define FP16_TO_INDEX_418F 2877
`define FP16_TO_INDEX_4190 2878
`define FP16_TO_INDEX_4191 2879
`define FP16_TO_INDEX_4192 2880
`define FP16_TO_INDEX_4193 2881
`define FP16_TO_INDEX_4194 2882
`define FP16_TO_INDEX_4195 2883
`define FP16_TO_INDEX_4196 2884
`define FP16_TO_INDEX_4197 2885
`define FP16_TO_INDEX_4198 2886
`define FP16_TO_INDEX_4199 2887
`define FP16_TO_INDEX_419A 2888
`define FP16_TO_INDEX_419B 2889
`define FP16_TO_INDEX_419C 2890
`define FP16_TO_INDEX_419D 2891
`define FP16_TO_INDEX_419E 2892
`define FP16_TO_INDEX_419F 2893
`define FP16_TO_INDEX_41A0 2894
`define FP16_TO_INDEX_41A1 2895
`define FP16_TO_INDEX_41A2 2896
`define FP16_TO_INDEX_41A3 2897
`define FP16_TO_INDEX_41A4 2898
`define FP16_TO_INDEX_41A5 2899
`define FP16_TO_INDEX_41A7 2900
`define FP16_TO_INDEX_41A8 2901
`define FP16_TO_INDEX_41A9 2902
`define FP16_TO_INDEX_41AA 2903
`define FP16_TO_INDEX_41AB 2904
`define FP16_TO_INDEX_41AC 2905
`define FP16_TO_INDEX_41AD 2906
`define FP16_TO_INDEX_41AE 2907
`define FP16_TO_INDEX_41AF 2908
`define FP16_TO_INDEX_41B0 2909
`define FP16_TO_INDEX_41B1 2910
`define FP16_TO_INDEX_41B2 2911
`define FP16_TO_INDEX_41B3 2912
`define FP16_TO_INDEX_41B4 2913
`define FP16_TO_INDEX_41B5 2914
`define FP16_TO_INDEX_41B6 2915
`define FP16_TO_INDEX_41B7 2916
`define FP16_TO_INDEX_41B8 2917
`define FP16_TO_INDEX_41B9 2918
`define FP16_TO_INDEX_41BA 2919
`define FP16_TO_INDEX_41BB 2920
`define FP16_TO_INDEX_41BC 2921
`define FP16_TO_INDEX_41BD 2922
`define FP16_TO_INDEX_41BE 2923
`define FP16_TO_INDEX_41BF 2924
`define FP16_TO_INDEX_41C0 2925
`define FP16_TO_INDEX_41C1 2926
`define FP16_TO_INDEX_41C2 2927
`define FP16_TO_INDEX_41C3 2928
`define FP16_TO_INDEX_41C4 2929
`define FP16_TO_INDEX_41C5 2930
`define FP16_TO_INDEX_41C6 2931
`define FP16_TO_INDEX_41C7 2932
`define FP16_TO_INDEX_41C8 2933
`define FP16_TO_INDEX_41C9 2934
`define FP16_TO_INDEX_41CB 2935
`define FP16_TO_INDEX_41CC 2936
`define FP16_TO_INDEX_41CD 2937
`define FP16_TO_INDEX_41CE 2938
`define FP16_TO_INDEX_41CF 2939
`define FP16_TO_INDEX_41D0 2940
`define FP16_TO_INDEX_41D1 2941
`define FP16_TO_INDEX_41D2 2942
`define FP16_TO_INDEX_41D3 2943
`define FP16_TO_INDEX_41D4 2944
`define FP16_TO_INDEX_41D5 2945
`define FP16_TO_INDEX_41D6 2946
`define FP16_TO_INDEX_41D7 2947
`define FP16_TO_INDEX_41D8 2948
`define FP16_TO_INDEX_41D9 2949
`define FP16_TO_INDEX_41DA 2950
`define FP16_TO_INDEX_41DB 2951
`define FP16_TO_INDEX_41DC 2952
`define FP16_TO_INDEX_41DD 2953
`define FP16_TO_INDEX_41DE 2954
`define FP16_TO_INDEX_41DF 2955
`define FP16_TO_INDEX_41E0 2956
`define FP16_TO_INDEX_41E1 2957
`define FP16_TO_INDEX_41E2 2958
`define FP16_TO_INDEX_41E3 2959
`define FP16_TO_INDEX_41E4 2960
`define FP16_TO_INDEX_41E5 2961
`define FP16_TO_INDEX_41E6 2962
`define FP16_TO_INDEX_41E7 2963
`define FP16_TO_INDEX_41E8 2964
`define FP16_TO_INDEX_41E9 2965
`define FP16_TO_INDEX_41EA 2966
`define FP16_TO_INDEX_41EB 2967
`define FP16_TO_INDEX_41EC 2968
`define FP16_TO_INDEX_41ED 2969
`define FP16_TO_INDEX_41EF 2970
`define FP16_TO_INDEX_41F0 2971
`define FP16_TO_INDEX_41F1 2972
`define FP16_TO_INDEX_41F2 2973
`define FP16_TO_INDEX_41F3 2974
`define FP16_TO_INDEX_41F4 2975
`define FP16_TO_INDEX_41F5 2976
`define FP16_TO_INDEX_41F6 2977
`define FP16_TO_INDEX_41F7 2978
`define FP16_TO_INDEX_41F8 2979
`define FP16_TO_INDEX_41F9 2980
`define FP16_TO_INDEX_41FA 2981
`define FP16_TO_INDEX_41FB 2982
`define FP16_TO_INDEX_41FC 2983
`define FP16_TO_INDEX_41FD 2984
`define FP16_TO_INDEX_41FE 2985
`define FP16_TO_INDEX_41FF 2986
`define FP16_TO_INDEX_4200 2987
