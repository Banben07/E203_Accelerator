`define CUBE_LUT_SIZE 1024
`define CUBE_LUT_BITS 10
`define CUBE_LUT_C200 16'hCEC0
`define CUBE_LUT_C1FF 16'hCEBD
`define CUBE_LUT_C1FE 16'hCEB9
`define CUBE_LUT_C1FD 16'hCEB6
`define CUBE_LUT_C1FC 16'hCEB3
`define CUBE_LUT_C1FB 16'hCEAF
`define CUBE_LUT_C1FA 16'hCEAC
`define CUBE_LUT_C1F9 16'hCEA8
`define CUBE_LUT_C1F8 16'hCEA5
`define CUBE_LUT_C1F7 16'hCEA2
`define CUBE_LUT_C1F6 16'hCE9E
`define CUBE_LUT_C1F5 16'hCE9B
`define CUBE_LUT_C1F4 16'hCE98
`define CUBE_LUT_C1F3 16'hCE94
`define CUBE_LUT_C1F2 16'hCE91
`define CUBE_LUT_C1F1 16'hCE8E
`define CUBE_LUT_C1F0 16'hCE8B
`define CUBE_LUT_C1EF 16'hCE87
`define CUBE_LUT_C1EE 16'hCE84
`define CUBE_LUT_C1ED 16'hCE81
`define CUBE_LUT_C1EC 16'hCE7D
`define CUBE_LUT_C1EB 16'hCE7A
`define CUBE_LUT_C1EA 16'hCE77
`define CUBE_LUT_C1E9 16'hCE74
`define CUBE_LUT_C1E8 16'hCE70
`define CUBE_LUT_C1E7 16'hCE6D
`define CUBE_LUT_C1E6 16'hCE6A
`define CUBE_LUT_C1E5 16'hCE66
`define CUBE_LUT_C1E4 16'hCE63
`define CUBE_LUT_C1E3 16'hCE60
`define CUBE_LUT_C1E2 16'hCE5D
`define CUBE_LUT_C1E1 16'hCE59
`define CUBE_LUT_C1E0 16'hCE56
`define CUBE_LUT_C1DF 16'hCE53
`define CUBE_LUT_C1DE 16'hCE50
`define CUBE_LUT_C1DD 16'hCE4D
`define CUBE_LUT_C1DC 16'hCE49
`define CUBE_LUT_C1DB 16'hCE46
`define CUBE_LUT_C1DA 16'hCE43
`define CUBE_LUT_C1D9 16'hCE40
`define CUBE_LUT_C1D8 16'hCE3C
`define CUBE_LUT_C1D7 16'hCE39
`define CUBE_LUT_C1D6 16'hCE36
`define CUBE_LUT_C1D5 16'hCE33
`define CUBE_LUT_C1D4 16'hCE30
`define CUBE_LUT_C1D3 16'hCE2D
`define CUBE_LUT_C1D2 16'hCE29
`define CUBE_LUT_C1D1 16'hCE26
`define CUBE_LUT_C1D0 16'hCE23
`define CUBE_LUT_C1CF 16'hCE20
`define CUBE_LUT_C1CE 16'hCE1D
`define CUBE_LUT_C1CD 16'hCE1A
`define CUBE_LUT_C1CC 16'hCE16
`define CUBE_LUT_C1CB 16'hCE13
`define CUBE_LUT_C1CA 16'hCE10
`define CUBE_LUT_C1C9 16'hCE0D
`define CUBE_LUT_C1C8 16'hCE0A
`define CUBE_LUT_C1C7 16'hCE07
`define CUBE_LUT_C1C6 16'hCE04
`define CUBE_LUT_C1C5 16'hCE00
`define CUBE_LUT_C1C4 16'hCDFD
`define CUBE_LUT_C1C3 16'hCDFA
`define CUBE_LUT_C1C2 16'hCDF7
`define CUBE_LUT_C1C1 16'hCDF4
`define CUBE_LUT_C1C0 16'hCDF1
`define CUBE_LUT_C1BF 16'hCDEE
`define CUBE_LUT_C1BE 16'hCDEB
`define CUBE_LUT_C1BD 16'hCDE8
`define CUBE_LUT_C1BC 16'hCDE5
`define CUBE_LUT_C1BB 16'hCDE1
`define CUBE_LUT_C1BA 16'hCDDE
`define CUBE_LUT_C1B9 16'hCDDB
`define CUBE_LUT_C1B8 16'hCDD8
`define CUBE_LUT_C1B7 16'hCDD5
`define CUBE_LUT_C1B6 16'hCDD2
`define CUBE_LUT_C1B5 16'hCDCF
`define CUBE_LUT_C1B4 16'hCDCC
`define CUBE_LUT_C1B3 16'hCDC9
`define CUBE_LUT_C1B2 16'hCDC6
`define CUBE_LUT_C1B1 16'hCDC3
`define CUBE_LUT_C1B0 16'hCDC0
`define CUBE_LUT_C1AF 16'hCDBD
`define CUBE_LUT_C1AE 16'hCDBA
`define CUBE_LUT_C1AD 16'hCDB7
`define CUBE_LUT_C1AC 16'hCDB4
`define CUBE_LUT_C1AB 16'hCDB1
`define CUBE_LUT_C1AA 16'hCDAE
`define CUBE_LUT_C1A9 16'hCDAB
`define CUBE_LUT_C1A8 16'hCDA8
`define CUBE_LUT_C1A7 16'hCDA5
`define CUBE_LUT_C1A6 16'hCDA2
`define CUBE_LUT_C1A5 16'hCD9F
`define CUBE_LUT_C1A4 16'hCD9C
`define CUBE_LUT_C1A3 16'hCD99
`define CUBE_LUT_C1A2 16'hCD96
`define CUBE_LUT_C1A1 16'hCD93
`define CUBE_LUT_C1A0 16'hCD90
`define CUBE_LUT_C19F 16'hCD8D
`define CUBE_LUT_C19E 16'hCD8A
`define CUBE_LUT_C19D 16'hCD87
`define CUBE_LUT_C19C 16'hCD84
`define CUBE_LUT_C19B 16'hCD81
`define CUBE_LUT_C19A 16'hCD7E
`define CUBE_LUT_C199 16'hCD7B
`define CUBE_LUT_C198 16'hCD78
`define CUBE_LUT_C197 16'hCD75
`define CUBE_LUT_C196 16'hCD72
`define CUBE_LUT_C195 16'hCD6F
`define CUBE_LUT_C194 16'hCD6D
`define CUBE_LUT_C193 16'hCD6A
`define CUBE_LUT_C192 16'hCD67
`define CUBE_LUT_C191 16'hCD64
`define CUBE_LUT_C190 16'hCD61
`define CUBE_LUT_C18F 16'hCD5E
`define CUBE_LUT_C18E 16'hCD5B
`define CUBE_LUT_C18D 16'hCD58
`define CUBE_LUT_C18C 16'hCD55
`define CUBE_LUT_C18B 16'hCD52
`define CUBE_LUT_C18A 16'hCD50
`define CUBE_LUT_C189 16'hCD4D
`define CUBE_LUT_C188 16'hCD4A
`define CUBE_LUT_C187 16'hCD47
`define CUBE_LUT_C186 16'hCD44
`define CUBE_LUT_C185 16'hCD41
`define CUBE_LUT_C184 16'hCD3E
`define CUBE_LUT_C183 16'hCD3C
`define CUBE_LUT_C182 16'hCD39
`define CUBE_LUT_C181 16'hCD36
`define CUBE_LUT_C180 16'hCD33
`define CUBE_LUT_C17F 16'hCD30
`define CUBE_LUT_C17E 16'hCD2D
`define CUBE_LUT_C17D 16'hCD2B
`define CUBE_LUT_C17C 16'hCD28
`define CUBE_LUT_C17B 16'hCD25
`define CUBE_LUT_C17A 16'hCD22
`define CUBE_LUT_C179 16'hCD1F
`define CUBE_LUT_C178 16'hCD1C
`define CUBE_LUT_C177 16'hCD1A
`define CUBE_LUT_C176 16'hCD17
`define CUBE_LUT_C175 16'hCD14
`define CUBE_LUT_C174 16'hCD11
`define CUBE_LUT_C173 16'hCD0E
`define CUBE_LUT_C172 16'hCD0C
`define CUBE_LUT_C171 16'hCD09
`define CUBE_LUT_C170 16'hCD06
`define CUBE_LUT_C16F 16'hCD03
`define CUBE_LUT_C16E 16'hCD01
`define CUBE_LUT_C16D 16'hCCFE
`define CUBE_LUT_C16C 16'hCCFB
`define CUBE_LUT_C16B 16'hCCF8
`define CUBE_LUT_C16A 16'hCCF6
`define CUBE_LUT_C169 16'hCCF3
`define CUBE_LUT_C168 16'hCCF0
`define CUBE_LUT_C167 16'hCCED
`define CUBE_LUT_C166 16'hCCEB
`define CUBE_LUT_C165 16'hCCE8
`define CUBE_LUT_C164 16'hCCE5
`define CUBE_LUT_C163 16'hCCE2
`define CUBE_LUT_C162 16'hCCE0
`define CUBE_LUT_C161 16'hCCDD
`define CUBE_LUT_C160 16'hCCDA
`define CUBE_LUT_C15F 16'hCCD8
`define CUBE_LUT_C15E 16'hCCD5
`define CUBE_LUT_C15D 16'hCCD2
`define CUBE_LUT_C15C 16'hCCCF
`define CUBE_LUT_C15B 16'hCCCD
`define CUBE_LUT_C15A 16'hCCCA
`define CUBE_LUT_C159 16'hCCC7
`define CUBE_LUT_C158 16'hCCC5
`define CUBE_LUT_C157 16'hCCC2
`define CUBE_LUT_C156 16'hCCBF
`define CUBE_LUT_C155 16'hCCBD
`define CUBE_LUT_C154 16'hCCBA
`define CUBE_LUT_C153 16'hCCB7
`define CUBE_LUT_C152 16'hCCB5
`define CUBE_LUT_C151 16'hCCB2
`define CUBE_LUT_C150 16'hCCAF
`define CUBE_LUT_C14F 16'hCCAD
`define CUBE_LUT_C14E 16'hCCAA
`define CUBE_LUT_C14D 16'hCCA8
`define CUBE_LUT_C14C 16'hCCA5
`define CUBE_LUT_C14B 16'hCCA2
`define CUBE_LUT_C14A 16'hCCA0
`define CUBE_LUT_C149 16'hCC9D
`define CUBE_LUT_C148 16'hCC9A
`define CUBE_LUT_C147 16'hCC98
`define CUBE_LUT_C146 16'hCC95
`define CUBE_LUT_C145 16'hCC93
`define CUBE_LUT_C144 16'hCC90
`define CUBE_LUT_C143 16'hCC8D
`define CUBE_LUT_C142 16'hCC8B
`define CUBE_LUT_C141 16'hCC88
`define CUBE_LUT_C140 16'hCC86
`define CUBE_LUT_C13F 16'hCC83
`define CUBE_LUT_C13E 16'hCC80
`define CUBE_LUT_C13D 16'hCC7E
`define CUBE_LUT_C13C 16'hCC7B
`define CUBE_LUT_C13B 16'hCC79
`define CUBE_LUT_C13A 16'hCC76
`define CUBE_LUT_C139 16'hCC74
`define CUBE_LUT_C138 16'hCC71
`define CUBE_LUT_C137 16'hCC6F
`define CUBE_LUT_C136 16'hCC6C
`define CUBE_LUT_C135 16'hCC69
`define CUBE_LUT_C134 16'hCC67
`define CUBE_LUT_C133 16'hCC64
`define CUBE_LUT_C132 16'hCC62
`define CUBE_LUT_C131 16'hCC5F
`define CUBE_LUT_C130 16'hCC5D
`define CUBE_LUT_C12F 16'hCC5A
`define CUBE_LUT_C12E 16'hCC58
`define CUBE_LUT_C12D 16'hCC55
`define CUBE_LUT_C12C 16'hCC53
`define CUBE_LUT_C12B 16'hCC50
`define CUBE_LUT_C12A 16'hCC4E
`define CUBE_LUT_C129 16'hCC4B
`define CUBE_LUT_C128 16'hCC49
`define CUBE_LUT_C127 16'hCC46
`define CUBE_LUT_C126 16'hCC44
`define CUBE_LUT_C125 16'hCC41
`define CUBE_LUT_C124 16'hCC3F
`define CUBE_LUT_C123 16'hCC3C
`define CUBE_LUT_C122 16'hCC3A
`define CUBE_LUT_C121 16'hCC37
`define CUBE_LUT_C120 16'hCC35
`define CUBE_LUT_C11F 16'hCC32
`define CUBE_LUT_C11E 16'hCC30
`define CUBE_LUT_C11D 16'hCC2E
`define CUBE_LUT_C11C 16'hCC2B
`define CUBE_LUT_C11B 16'hCC29
`define CUBE_LUT_C11A 16'hCC26
`define CUBE_LUT_C119 16'hCC24
`define CUBE_LUT_C118 16'hCC21
`define CUBE_LUT_C117 16'hCC1F
`define CUBE_LUT_C116 16'hCC1C
`define CUBE_LUT_C115 16'hCC1A
`define CUBE_LUT_C114 16'hCC18
`define CUBE_LUT_C113 16'hCC15
`define CUBE_LUT_C112 16'hCC13
`define CUBE_LUT_C111 16'hCC10
`define CUBE_LUT_C110 16'hCC0E
`define CUBE_LUT_C10F 16'hCC0C
`define CUBE_LUT_C10E 16'hCC09
`define CUBE_LUT_C10D 16'hCC07
`define CUBE_LUT_C10C 16'hCC04
`define CUBE_LUT_C10B 16'hCC02
`define CUBE_LUT_C10A 16'hCBFF
`define CUBE_LUT_C109 16'hCBFA
`define CUBE_LUT_C108 16'hCBF6
`define CUBE_LUT_C107 16'hCBF1
`define CUBE_LUT_C106 16'hCBEC
`define CUBE_LUT_C105 16'hCBE8
`define CUBE_LUT_C104 16'hCBE3
`define CUBE_LUT_C103 16'hCBDE
`define CUBE_LUT_C102 16'hCBD9
`define CUBE_LUT_C101 16'hCBD5
`define CUBE_LUT_C100 16'hCBD0
`define CUBE_LUT_C0FF 16'hCBCB
`define CUBE_LUT_C0FE 16'hCBC7
`define CUBE_LUT_C0FD 16'hCBC2
`define CUBE_LUT_C0FC 16'hCBBD
`define CUBE_LUT_C0FB 16'hCBB9
`define CUBE_LUT_C0FA 16'hCBB4
`define CUBE_LUT_C0F9 16'hCBAF
`define CUBE_LUT_C0F8 16'hCBAB
`define CUBE_LUT_C0F7 16'hCBA6
`define CUBE_LUT_C0F6 16'hCBA1
`define CUBE_LUT_C0F5 16'hCB9D
`define CUBE_LUT_C0F4 16'hCB98
`define CUBE_LUT_C0F3 16'hCB94
`define CUBE_LUT_C0F2 16'hCB8F
`define CUBE_LUT_C0F1 16'hCB8B
`define CUBE_LUT_C0F0 16'hCB86
`define CUBE_LUT_C0EF 16'hCB81
`define CUBE_LUT_C0EE 16'hCB7D
`define CUBE_LUT_C0ED 16'hCB78
`define CUBE_LUT_C0EC 16'hCB74
`define CUBE_LUT_C0EB 16'hCB6F
`define CUBE_LUT_C0EA 16'hCB6B
`define CUBE_LUT_C0E9 16'hCB66
`define CUBE_LUT_C0E8 16'hCB62
`define CUBE_LUT_C0E7 16'hCB5D
`define CUBE_LUT_C0E6 16'hCB59
`define CUBE_LUT_C0E5 16'hCB54
`define CUBE_LUT_C0E4 16'hCB50
`define CUBE_LUT_C0E3 16'hCB4B
`define CUBE_LUT_C0E2 16'hCB47
`define CUBE_LUT_C0E1 16'hCB42
`define CUBE_LUT_C0E0 16'hCB3E
`define CUBE_LUT_C0DF 16'hCB39
`define CUBE_LUT_C0DE 16'hCB35
`define CUBE_LUT_C0DD 16'hCB30
`define CUBE_LUT_C0DC 16'hCB2C
`define CUBE_LUT_C0DB 16'hCB28
`define CUBE_LUT_C0DA 16'hCB23
`define CUBE_LUT_C0D9 16'hCB1F
`define CUBE_LUT_C0D8 16'hCB1A
`define CUBE_LUT_C0D7 16'hCB16
`define CUBE_LUT_C0D6 16'hCB12
`define CUBE_LUT_C0D5 16'hCB0D
`define CUBE_LUT_C0D4 16'hCB09
`define CUBE_LUT_C0D3 16'hCB04
`define CUBE_LUT_C0D2 16'hCB00
`define CUBE_LUT_C0D1 16'hCAFC
`define CUBE_LUT_C0D0 16'hCAF7
`define CUBE_LUT_C0CF 16'hCAF3
`define CUBE_LUT_C0CE 16'hCAEF
`define CUBE_LUT_C0CD 16'hCAEA
`define CUBE_LUT_C0CC 16'hCAE6
`define CUBE_LUT_C0CB 16'hCAE2
`define CUBE_LUT_C0CA 16'hCADD
`define CUBE_LUT_C0C9 16'hCAD9
`define CUBE_LUT_C0C8 16'hCAD5
`define CUBE_LUT_C0C7 16'hCAD1
`define CUBE_LUT_C0C6 16'hCACC
`define CUBE_LUT_C0C5 16'hCAC8
`define CUBE_LUT_C0C4 16'hCAC4
`define CUBE_LUT_C0C3 16'hCABF
`define CUBE_LUT_C0C2 16'hCABB
`define CUBE_LUT_C0C1 16'hCAB7
`define CUBE_LUT_C0C0 16'hCAB3
`define CUBE_LUT_C0BF 16'hCAAF
`define CUBE_LUT_C0BE 16'hCAAA
`define CUBE_LUT_C0BD 16'hCAA6
`define CUBE_LUT_C0BC 16'hCAA2
`define CUBE_LUT_C0BB 16'hCA9E
`define CUBE_LUT_C0BA 16'hCA99
`define CUBE_LUT_C0B9 16'hCA95
`define CUBE_LUT_C0B8 16'hCA91
`define CUBE_LUT_C0B7 16'hCA8D
`define CUBE_LUT_C0B6 16'hCA89
`define CUBE_LUT_C0B5 16'hCA85
`define CUBE_LUT_C0B4 16'hCA80
`define CUBE_LUT_C0B3 16'hCA7C
`define CUBE_LUT_C0B2 16'hCA78
`define CUBE_LUT_C0B1 16'hCA74
`define CUBE_LUT_C0B0 16'hCA70
`define CUBE_LUT_C0AF 16'hCA6C
`define CUBE_LUT_C0AE 16'hCA68
`define CUBE_LUT_C0AD 16'hCA64
`define CUBE_LUT_C0AC 16'hCA60
`define CUBE_LUT_C0AB 16'hCA5B
`define CUBE_LUT_C0AA 16'hCA57
`define CUBE_LUT_C0A9 16'hCA53
`define CUBE_LUT_C0A8 16'hCA4F
`define CUBE_LUT_C0A7 16'hCA4B
`define CUBE_LUT_C0A6 16'hCA47
`define CUBE_LUT_C0A5 16'hCA43
`define CUBE_LUT_C0A4 16'hCA3F
`define CUBE_LUT_C0A3 16'hCA3B
`define CUBE_LUT_C0A2 16'hCA37
`define CUBE_LUT_C0A1 16'hCA33
`define CUBE_LUT_C0A0 16'hCA2F
`define CUBE_LUT_C09F 16'hCA2B
`define CUBE_LUT_C09E 16'hCA27
`define CUBE_LUT_C09D 16'hCA23
`define CUBE_LUT_C09C 16'hCA1F
`define CUBE_LUT_C09B 16'hCA1B
`define CUBE_LUT_C09A 16'hCA17
`define CUBE_LUT_C099 16'hCA13
`define CUBE_LUT_C098 16'hCA0F
`define CUBE_LUT_C097 16'hCA0B
`define CUBE_LUT_C096 16'hCA07
`define CUBE_LUT_C095 16'hCA03
`define CUBE_LUT_C094 16'hC9FF
`define CUBE_LUT_C093 16'hC9FB
`define CUBE_LUT_C092 16'hC9F7
`define CUBE_LUT_C091 16'hC9F4
`define CUBE_LUT_C090 16'hC9F0
`define CUBE_LUT_C08F 16'hC9EC
`define CUBE_LUT_C08E 16'hC9E8
`define CUBE_LUT_C08D 16'hC9E4
`define CUBE_LUT_C08C 16'hC9E0
`define CUBE_LUT_C08B 16'hC9DC
`define CUBE_LUT_C08A 16'hC9D8
`define CUBE_LUT_C089 16'hC9D4
`define CUBE_LUT_C088 16'hC9D1
`define CUBE_LUT_C087 16'hC9CD
`define CUBE_LUT_C086 16'hC9C9
`define CUBE_LUT_C085 16'hC9C5
`define CUBE_LUT_C084 16'hC9C1
`define CUBE_LUT_C083 16'hC9BD
`define CUBE_LUT_C082 16'hC9BA
`define CUBE_LUT_C081 16'hC9B6
`define CUBE_LUT_C080 16'hC9B2
`define CUBE_LUT_C07F 16'hC9AE
`define CUBE_LUT_C07E 16'hC9AA
`define CUBE_LUT_C07D 16'hC9A7
`define CUBE_LUT_C07C 16'hC9A3
`define CUBE_LUT_C07B 16'hC99F
`define CUBE_LUT_C07A 16'hC99B
`define CUBE_LUT_C079 16'hC998
`define CUBE_LUT_C078 16'hC994
`define CUBE_LUT_C077 16'hC990
`define CUBE_LUT_C076 16'hC98C
`define CUBE_LUT_C075 16'hC989
`define CUBE_LUT_C074 16'hC985
`define CUBE_LUT_C073 16'hC981
`define CUBE_LUT_C072 16'hC97D
`define CUBE_LUT_C071 16'hC97A
`define CUBE_LUT_C070 16'hC976
`define CUBE_LUT_C06F 16'hC972
`define CUBE_LUT_C06E 16'hC96F
`define CUBE_LUT_C06D 16'hC96B
`define CUBE_LUT_C06C 16'hC967
`define CUBE_LUT_C06B 16'hC964
`define CUBE_LUT_C06A 16'hC960
`define CUBE_LUT_C069 16'hC95C
`define CUBE_LUT_C068 16'hC959
`define CUBE_LUT_C067 16'hC955
`define CUBE_LUT_C066 16'hC951
`define CUBE_LUT_C065 16'hC94E
`define CUBE_LUT_C064 16'hC94A
`define CUBE_LUT_C063 16'hC947
`define CUBE_LUT_C062 16'hC943
`define CUBE_LUT_C061 16'hC93F
`define CUBE_LUT_C060 16'hC93C
`define CUBE_LUT_C05F 16'hC938
`define CUBE_LUT_C05E 16'hC935
`define CUBE_LUT_C05D 16'hC931
`define CUBE_LUT_C05C 16'hC92E
`define CUBE_LUT_C05B 16'hC92A
`define CUBE_LUT_C05A 16'hC926
`define CUBE_LUT_C059 16'hC923
`define CUBE_LUT_C058 16'hC91F
`define CUBE_LUT_C057 16'hC91C
`define CUBE_LUT_C056 16'hC918
`define CUBE_LUT_C055 16'hC915
`define CUBE_LUT_C054 16'hC911
`define CUBE_LUT_C053 16'hC90E
`define CUBE_LUT_C052 16'hC90A
`define CUBE_LUT_C051 16'hC907
`define CUBE_LUT_C050 16'hC903
`define CUBE_LUT_C04F 16'hC900
`define CUBE_LUT_C04E 16'hC8FC
`define CUBE_LUT_C04D 16'hC8F9
`define CUBE_LUT_C04C 16'hC8F5
`define CUBE_LUT_C04B 16'hC8F2
`define CUBE_LUT_C04A 16'hC8EE
`define CUBE_LUT_C049 16'hC8EB
`define CUBE_LUT_C048 16'hC8E8
`define CUBE_LUT_C047 16'hC8E4
`define CUBE_LUT_C046 16'hC8E1
`define CUBE_LUT_C045 16'hC8DD
`define CUBE_LUT_C044 16'hC8DA
`define CUBE_LUT_C043 16'hC8D6
`define CUBE_LUT_C042 16'hC8D3
`define CUBE_LUT_C041 16'hC8D0
`define CUBE_LUT_C040 16'hC8CC
`define CUBE_LUT_C03F 16'hC8C9
`define CUBE_LUT_C03E 16'hC8C5
`define CUBE_LUT_C03D 16'hC8C2
`define CUBE_LUT_C03C 16'hC8BF
`define CUBE_LUT_C03B 16'hC8BB
`define CUBE_LUT_C03A 16'hC8B8
`define CUBE_LUT_C039 16'hC8B5
`define CUBE_LUT_C038 16'hC8B1
`define CUBE_LUT_C037 16'hC8AE
`define CUBE_LUT_C036 16'hC8AB
`define CUBE_LUT_C035 16'hC8A7
`define CUBE_LUT_C034 16'hC8A4
`define CUBE_LUT_C033 16'hC8A1
`define CUBE_LUT_C032 16'hC89D
`define CUBE_LUT_C031 16'hC89A
`define CUBE_LUT_C030 16'hC897
`define CUBE_LUT_C02F 16'hC894
`define CUBE_LUT_C02E 16'hC890
`define CUBE_LUT_C02D 16'hC88D
`define CUBE_LUT_C02C 16'hC88A
`define CUBE_LUT_C02B 16'hC886
`define CUBE_LUT_C02A 16'hC883
`define CUBE_LUT_C029 16'hC880
`define CUBE_LUT_C028 16'hC87D
`define CUBE_LUT_C027 16'hC87A
`define CUBE_LUT_C026 16'hC876
`define CUBE_LUT_C025 16'hC873
`define CUBE_LUT_C024 16'hC870
`define CUBE_LUT_C023 16'hC86D
`define CUBE_LUT_C022 16'hC869
`define CUBE_LUT_C021 16'hC866
`define CUBE_LUT_C020 16'hC863
`define CUBE_LUT_C01F 16'hC860
`define CUBE_LUT_C01E 16'hC85D
`define CUBE_LUT_C01D 16'hC859
`define CUBE_LUT_C01C 16'hC856
`define CUBE_LUT_C01B 16'hC853
`define CUBE_LUT_C01A 16'hC850
`define CUBE_LUT_C019 16'hC84D
`define CUBE_LUT_C018 16'hC84A
`define CUBE_LUT_C017 16'hC847
`define CUBE_LUT_C016 16'hC843
`define CUBE_LUT_C015 16'hC840
`define CUBE_LUT_C014 16'hC83D
`define CUBE_LUT_C013 16'hC83A
`define CUBE_LUT_C012 16'hC837
`define CUBE_LUT_C011 16'hC834
`define CUBE_LUT_C010 16'hC831
`define CUBE_LUT_C00F 16'hC82E
`define CUBE_LUT_C00E 16'hC82B
`define CUBE_LUT_C00D 16'hC827
`define CUBE_LUT_C00C 16'hC824
`define CUBE_LUT_C00B 16'hC821
`define CUBE_LUT_C00A 16'hC81E
`define CUBE_LUT_C009 16'hC81B
`define CUBE_LUT_C008 16'hC818
`define CUBE_LUT_C007 16'hC815
`define CUBE_LUT_C006 16'hC812
`define CUBE_LUT_C005 16'hC80F
`define CUBE_LUT_C004 16'hC80C
`define CUBE_LUT_C003 16'hC809
`define CUBE_LUT_C002 16'hC806
`define CUBE_LUT_C001 16'hC803
`define CUBE_LUT_C000 16'hC800
`define CUBE_LUT_BFFF 16'hC7FD
`define CUBE_LUT_BFFE 16'hC7FA
`define CUBE_LUT_BFFD 16'hC7F7
`define CUBE_LUT_BFFC 16'hC7F4
`define CUBE_LUT_BFFB 16'hC7F1
`define CUBE_LUT_BFFA 16'hC7EE
`define CUBE_LUT_BFF9 16'hC7EB
`define CUBE_LUT_BFF8 16'hC7E8
`define CUBE_LUT_BFF7 16'hC7E5
`define CUBE_LUT_BFF6 16'hC7E2
`define CUBE_LUT_BFF5 16'hC7DF
`define CUBE_LUT_BFF4 16'hC7DC
`define CUBE_LUT_BFF3 16'hC7D9
`define CUBE_LUT_BFF2 16'hC7D6
`define CUBE_LUT_BFF1 16'hC7D3
`define CUBE_LUT_BFF0 16'hC7D0
`define CUBE_LUT_BFEF 16'hC7CD
`define CUBE_LUT_BFEE 16'hC7CA
`define CUBE_LUT_BFED 16'hC7C8
`define CUBE_LUT_BFEC 16'hC7C5
`define CUBE_LUT_BFEB 16'hC7C2
`define CUBE_LUT_BFEA 16'hC7BF
`define CUBE_LUT_BFE9 16'hC7BC
`define CUBE_LUT_BFE8 16'hC7B9
`define CUBE_LUT_BFE7 16'hC7B6
`define CUBE_LUT_BFE6 16'hC7B3
`define CUBE_LUT_BFE5 16'hC7B0
`define CUBE_LUT_BFE4 16'hC7AD
`define CUBE_LUT_BFE3 16'hC7AA
`define CUBE_LUT_BFE2 16'hC7A7
`define CUBE_LUT_BFE1 16'hC7A4
`define CUBE_LUT_BFE0 16'hC7A1
`define CUBE_LUT_BFDF 16'hC79F
`define CUBE_LUT_BFDE 16'hC79C
`define CUBE_LUT_BFDD 16'hC799
`define CUBE_LUT_BFDC 16'hC796
`define CUBE_LUT_BFDB 16'hC793
`define CUBE_LUT_BFDA 16'hC790
`define CUBE_LUT_BFD9 16'hC78D
`define CUBE_LUT_BFD8 16'hC78A
`define CUBE_LUT_BFD7 16'hC787
`define CUBE_LUT_BFD6 16'hC785
`define CUBE_LUT_BFD5 16'hC782
`define CUBE_LUT_BFD4 16'hC77F
`define CUBE_LUT_BFD3 16'hC77C
`define CUBE_LUT_BFD2 16'hC779
`define CUBE_LUT_BFD1 16'hC776
`define CUBE_LUT_BFD0 16'hC773
`define CUBE_LUT_BFCF 16'hC770
`define CUBE_LUT_BFCE 16'hC76E
`define CUBE_LUT_BFCD 16'hC76B
`define CUBE_LUT_BFCC 16'hC768
`define CUBE_LUT_BFCB 16'hC765
`define CUBE_LUT_BFCA 16'hC762
`define CUBE_LUT_BFC9 16'hC75F
`define CUBE_LUT_BFC8 16'hC75D
`define CUBE_LUT_BFC7 16'hC75A
`define CUBE_LUT_BFC6 16'hC757
`define CUBE_LUT_BFC5 16'hC754
`define CUBE_LUT_BFC4 16'hC751
`define CUBE_LUT_BFC3 16'hC74E
`define CUBE_LUT_BFC2 16'hC74C
`define CUBE_LUT_BFC1 16'hC749
`define CUBE_LUT_BFC0 16'hC746
`define CUBE_LUT_BFBF 16'hC743
`define CUBE_LUT_BFBE 16'hC740
`define CUBE_LUT_BFBD 16'hC73E
`define CUBE_LUT_BFBC 16'hC73B
`define CUBE_LUT_BFBB 16'hC738
`define CUBE_LUT_BFBA 16'hC735
`define CUBE_LUT_BFB9 16'hC732
`define CUBE_LUT_BFB8 16'hC730
`define CUBE_LUT_BFB7 16'hC72D
`define CUBE_LUT_BFB6 16'hC72A
`define CUBE_LUT_BFB5 16'hC727
`define CUBE_LUT_BFB4 16'hC724
`define CUBE_LUT_BFB3 16'hC722
`define CUBE_LUT_BFB2 16'hC71F
`define CUBE_LUT_BFB1 16'hC71C
`define CUBE_LUT_BFB0 16'hC719
`define CUBE_LUT_BFAF 16'hC716
`define CUBE_LUT_BFAE 16'hC714
`define CUBE_LUT_BFAD 16'hC711
`define CUBE_LUT_BFAC 16'hC70E
`define CUBE_LUT_BFAB 16'hC70B
`define CUBE_LUT_BFAA 16'hC709
`define CUBE_LUT_BFA9 16'hC706
`define CUBE_LUT_BFA8 16'hC703
`define CUBE_LUT_BFA7 16'hC700
`define CUBE_LUT_BFA6 16'hC6FE
`define CUBE_LUT_BFA5 16'hC6FB
`define CUBE_LUT_BFA4 16'hC6F8
`define CUBE_LUT_BFA3 16'hC6F5
`define CUBE_LUT_BFA2 16'hC6F3
`define CUBE_LUT_BFA1 16'hC6F0
`define CUBE_LUT_BFA0 16'hC6ED
`define CUBE_LUT_BF9F 16'hC6EB
`define CUBE_LUT_BF9E 16'hC6E8
`define CUBE_LUT_BF9D 16'hC6E5
`define CUBE_LUT_BF9C 16'hC6E2
`define CUBE_LUT_BF9B 16'hC6E0
`define CUBE_LUT_BF9A 16'hC6DD
`define CUBE_LUT_BF99 16'hC6DA
`define CUBE_LUT_BF98 16'hC6D8
`define CUBE_LUT_BF97 16'hC6D5
`define CUBE_LUT_BF96 16'hC6D2
`define CUBE_LUT_BF95 16'hC6CF
`define CUBE_LUT_BF94 16'hC6CD
`define CUBE_LUT_BF93 16'hC6CA
`define CUBE_LUT_BF92 16'hC6C7
`define CUBE_LUT_BF91 16'hC6C5
`define CUBE_LUT_BF90 16'hC6C2
`define CUBE_LUT_BF8F 16'hC6BF
`define CUBE_LUT_BF8E 16'hC6BD
`define CUBE_LUT_BF8D 16'hC6BA
`define CUBE_LUT_BF8C 16'hC6B7
`define CUBE_LUT_BF8B 16'hC6B5
`define CUBE_LUT_BF8A 16'hC6B2
`define CUBE_LUT_BF89 16'hC6AF
`define CUBE_LUT_BF88 16'hC6AD
`define CUBE_LUT_BF87 16'hC6AA
`define CUBE_LUT_BF86 16'hC6A7
`define CUBE_LUT_BF85 16'hC6A5
`define CUBE_LUT_BF84 16'hC6A2
`define CUBE_LUT_BF83 16'hC69F
`define CUBE_LUT_BF82 16'hC69D
`define CUBE_LUT_BF81 16'hC69A
`define CUBE_LUT_BF80 16'hC698
`define CUBE_LUT_BF7F 16'hC695
`define CUBE_LUT_BF7E 16'hC692
`define CUBE_LUT_BF7D 16'hC690
`define CUBE_LUT_BF7C 16'hC68D
`define CUBE_LUT_BF7B 16'hC68A
`define CUBE_LUT_BF7A 16'hC688
`define CUBE_LUT_BF79 16'hC685
`define CUBE_LUT_BF78 16'hC682
`define CUBE_LUT_BF77 16'hC680
`define CUBE_LUT_BF76 16'hC67D
`define CUBE_LUT_BF75 16'hC67B
`define CUBE_LUT_BF74 16'hC678
`define CUBE_LUT_BF73 16'hC675
`define CUBE_LUT_BF72 16'hC673
`define CUBE_LUT_BF71 16'hC670
`define CUBE_LUT_BF70 16'hC66E
`define CUBE_LUT_BF6F 16'hC66B
`define CUBE_LUT_BF6E 16'hC668
`define CUBE_LUT_BF6D 16'hC666
`define CUBE_LUT_BF6C 16'hC663
`define CUBE_LUT_BF6B 16'hC661
`define CUBE_LUT_BF6A 16'hC65E
`define CUBE_LUT_BF69 16'hC65C
`define CUBE_LUT_BF68 16'hC659
`define CUBE_LUT_BF67 16'hC656
`define CUBE_LUT_BF66 16'hC654
`define CUBE_LUT_BF65 16'hC651
`define CUBE_LUT_BF64 16'hC64F
`define CUBE_LUT_BF63 16'hC64C
`define CUBE_LUT_BF62 16'hC64A
`define CUBE_LUT_BF61 16'hC647
`define CUBE_LUT_BF60 16'hC645
`define CUBE_LUT_BF5F 16'hC642
`define CUBE_LUT_BF5E 16'hC63F
`define CUBE_LUT_BF5D 16'hC63D
`define CUBE_LUT_BF5C 16'hC63A
`define CUBE_LUT_BF5B 16'hC638
`define CUBE_LUT_BF5A 16'hC635
`define CUBE_LUT_BF59 16'hC633
`define CUBE_LUT_BF58 16'hC630
`define CUBE_LUT_BF57 16'hC62E
`define CUBE_LUT_BF56 16'hC62B
`define CUBE_LUT_BF55 16'hC629
`define CUBE_LUT_BF54 16'hC626
`define CUBE_LUT_BF53 16'hC624
`define CUBE_LUT_BF52 16'hC621
`define CUBE_LUT_BF51 16'hC61F
`define CUBE_LUT_BF50 16'hC61C
`define CUBE_LUT_BF4F 16'hC61A
`define CUBE_LUT_BF4E 16'hC617
`define CUBE_LUT_BF4D 16'hC615
`define CUBE_LUT_BF4C 16'hC612
`define CUBE_LUT_BF4B 16'hC610
`define CUBE_LUT_BF4A 16'hC60D
`define CUBE_LUT_BF49 16'hC60B
`define CUBE_LUT_BF48 16'hC608
`define CUBE_LUT_BF47 16'hC606
`define CUBE_LUT_BF46 16'hC603
`define CUBE_LUT_BF45 16'hC601
`define CUBE_LUT_BF44 16'hC5FE
`define CUBE_LUT_BF43 16'hC5FC
`define CUBE_LUT_BF42 16'hC5F9
`define CUBE_LUT_BF41 16'hC5F7
`define CUBE_LUT_BF40 16'hC5F4
`define CUBE_LUT_BF3F 16'hC5F2
`define CUBE_LUT_BF3E 16'hC5EF
`define CUBE_LUT_BF3D 16'hC5ED
`define CUBE_LUT_BF3C 16'hC5EA
`define CUBE_LUT_BF3B 16'hC5E8
`define CUBE_LUT_BF3A 16'hC5E6
`define CUBE_LUT_BF39 16'hC5E3
`define CUBE_LUT_BF38 16'hC5E1
`define CUBE_LUT_BF37 16'hC5DE
`define CUBE_LUT_BF36 16'hC5DC
`define CUBE_LUT_BF35 16'hC5D9
`define CUBE_LUT_BF34 16'hC5D7
`define CUBE_LUT_BF33 16'hC5D5
`define CUBE_LUT_BF32 16'hC5D2
`define CUBE_LUT_BF31 16'hC5D0
`define CUBE_LUT_BF30 16'hC5CD
`define CUBE_LUT_BF2F 16'hC5CB
`define CUBE_LUT_BF2E 16'hC5C8
`define CUBE_LUT_BF2D 16'hC5C6
`define CUBE_LUT_BF2C 16'hC5C4
`define CUBE_LUT_BF2B 16'hC5C1
`define CUBE_LUT_BF2A 16'hC5BF
`define CUBE_LUT_BF29 16'hC5BC
`define CUBE_LUT_BF28 16'hC5BA
`define CUBE_LUT_BF27 16'hC5B8
`define CUBE_LUT_BF26 16'hC5B5
`define CUBE_LUT_BF25 16'hC5B3
`define CUBE_LUT_BF24 16'hC5B0
`define CUBE_LUT_BF23 16'hC5AE
`define CUBE_LUT_BF22 16'hC5AC
`define CUBE_LUT_BF21 16'hC5A9
`define CUBE_LUT_BF20 16'hC5A7
`define CUBE_LUT_BF1F 16'hC5A4
`define CUBE_LUT_BF1E 16'hC5A2
`define CUBE_LUT_BF1D 16'hC5A0
`define CUBE_LUT_BF1C 16'hC59D
`define CUBE_LUT_BF1B 16'hC59B
`define CUBE_LUT_BF1A 16'hC599
`define CUBE_LUT_BF19 16'hC596
`define CUBE_LUT_BF18 16'hC594
`define CUBE_LUT_BF17 16'hC592
`define CUBE_LUT_BF16 16'hC58F
`define CUBE_LUT_BF15 16'hC58D
`define CUBE_LUT_BF14 16'hC58A
`define CUBE_LUT_BF13 16'hC588
`define CUBE_LUT_BF12 16'hC586
`define CUBE_LUT_BF11 16'hC583
`define CUBE_LUT_BF10 16'hC581
`define CUBE_LUT_BF0F 16'hC57F
`define CUBE_LUT_BF0E 16'hC57C
`define CUBE_LUT_BF0D 16'hC57A
`define CUBE_LUT_BF0C 16'hC578
`define CUBE_LUT_BF0B 16'hC575
`define CUBE_LUT_BF0A 16'hC573
`define CUBE_LUT_BF09 16'hC571
`define CUBE_LUT_BF08 16'hC56E
`define CUBE_LUT_BF07 16'hC56C
`define CUBE_LUT_BF06 16'hC56A
`define CUBE_LUT_BF05 16'hC568
`define CUBE_LUT_BF04 16'hC565
`define CUBE_LUT_BF03 16'hC563
`define CUBE_LUT_BF02 16'hC561
`define CUBE_LUT_BF01 16'hC55E
`define CUBE_LUT_BF00 16'hC55C
`define CUBE_LUT_BEFF 16'hC55A
`define CUBE_LUT_BEFE 16'hC557
`define CUBE_LUT_BEFD 16'hC555
`define CUBE_LUT_BEFC 16'hC553
`define CUBE_LUT_BEFB 16'hC551
`define CUBE_LUT_BEFA 16'hC54E
`define CUBE_LUT_BEF9 16'hC54C
`define CUBE_LUT_BEF8 16'hC54A
`define CUBE_LUT_BEF7 16'hC547
`define CUBE_LUT_BEF6 16'hC545
`define CUBE_LUT_BEF5 16'hC543
`define CUBE_LUT_BEF4 16'hC541
`define CUBE_LUT_BEF3 16'hC53E
`define CUBE_LUT_BEF2 16'hC53C
`define CUBE_LUT_BEF1 16'hC53A
`define CUBE_LUT_BEF0 16'hC538
`define CUBE_LUT_BEEF 16'hC535
`define CUBE_LUT_BEEE 16'hC533
`define CUBE_LUT_BEED 16'hC531
`define CUBE_LUT_BEEC 16'hC52F
`define CUBE_LUT_BEEB 16'hC52C
`define CUBE_LUT_BEEA 16'hC52A
`define CUBE_LUT_BEE9 16'hC528
`define CUBE_LUT_BEE8 16'hC526
`define CUBE_LUT_BEE7 16'hC523
`define CUBE_LUT_BEE6 16'hC521
`define CUBE_LUT_BEE5 16'hC51F
`define CUBE_LUT_BEE4 16'hC51D
`define CUBE_LUT_BEE3 16'hC51A
`define CUBE_LUT_BEE2 16'hC518
`define CUBE_LUT_BEE1 16'hC516
`define CUBE_LUT_BEE0 16'hC514
`define CUBE_LUT_BEDF 16'hC512
`define CUBE_LUT_BEDE 16'hC50F
`define CUBE_LUT_BEDD 16'hC50D
`define CUBE_LUT_BEDC 16'hC50B
`define CUBE_LUT_BEDB 16'hC509
`define CUBE_LUT_BEDA 16'hC507
`define CUBE_LUT_BED9 16'hC504
`define CUBE_LUT_BED8 16'hC502
`define CUBE_LUT_BED7 16'hC500
`define CUBE_LUT_BED6 16'hC4FE
`define CUBE_LUT_BED5 16'hC4FC
`define CUBE_LUT_BED4 16'hC4F9
`define CUBE_LUT_BED3 16'hC4F7
`define CUBE_LUT_BED2 16'hC4F5
`define CUBE_LUT_BED1 16'hC4F3
`define CUBE_LUT_BED0 16'hC4F1
`define CUBE_LUT_BECF 16'hC4EF
`define CUBE_LUT_BECE 16'hC4EC
`define CUBE_LUT_BECD 16'hC4EA
`define CUBE_LUT_BECC 16'hC4E8
`define CUBE_LUT_BECB 16'hC4E6
`define CUBE_LUT_BECA 16'hC4E4
`define CUBE_LUT_BEC9 16'hC4E2
`define CUBE_LUT_BEC8 16'hC4DF
`define CUBE_LUT_BEC7 16'hC4DD
`define CUBE_LUT_BEC6 16'hC4DB
`define CUBE_LUT_BEC5 16'hC4D9
`define CUBE_LUT_BEC4 16'hC4D7
`define CUBE_LUT_BEC3 16'hC4D5
`define CUBE_LUT_BEC2 16'hC4D2
`define CUBE_LUT_BEC1 16'hC4D0
`define CUBE_LUT_BEC0 16'hC4CE
`define CUBE_LUT_BEBF 16'hC4CC
`define CUBE_LUT_BEBE 16'hC4CA
`define CUBE_LUT_BEBD 16'hC4C8
`define CUBE_LUT_BEBC 16'hC4C6
`define CUBE_LUT_BEBB 16'hC4C4
`define CUBE_LUT_BEBA 16'hC4C1
`define CUBE_LUT_BEB9 16'hC4BF
`define CUBE_LUT_BEB8 16'hC4BD
`define CUBE_LUT_BEB7 16'hC4BB
`define CUBE_LUT_BEB6 16'hC4B9
`define CUBE_LUT_BEB5 16'hC4B7
`define CUBE_LUT_BEB4 16'hC4B5
`define CUBE_LUT_BEB3 16'hC4B3
`define CUBE_LUT_BEB2 16'hC4B1
`define CUBE_LUT_BEB1 16'hC4AE
`define CUBE_LUT_BEB0 16'hC4AC
`define CUBE_LUT_BEAF 16'hC4AA
`define CUBE_LUT_BEAE 16'hC4A8
`define CUBE_LUT_BEAD 16'hC4A6
`define CUBE_LUT_BEAC 16'hC4A4
`define CUBE_LUT_BEAB 16'hC4A2
`define CUBE_LUT_BEAA 16'hC4A0
`define CUBE_LUT_BEA9 16'hC49E
`define CUBE_LUT_BEA8 16'hC49C
`define CUBE_LUT_BEA7 16'hC49A
`define CUBE_LUT_BEA6 16'hC497
`define CUBE_LUT_BEA5 16'hC495
`define CUBE_LUT_BEA4 16'hC493
`define CUBE_LUT_BEA3 16'hC491
`define CUBE_LUT_BEA2 16'hC48F
`define CUBE_LUT_BEA1 16'hC48D
`define CUBE_LUT_BEA0 16'hC48B
`define CUBE_LUT_BE9F 16'hC489
`define CUBE_LUT_BE9E 16'hC487
`define CUBE_LUT_BE9D 16'hC485
`define CUBE_LUT_BE9C 16'hC483
`define CUBE_LUT_BE9B 16'hC481
`define CUBE_LUT_BE9A 16'hC47F
`define CUBE_LUT_BE99 16'hC47D
`define CUBE_LUT_BE98 16'hC47B
`define CUBE_LUT_BE97 16'hC479
`define CUBE_LUT_BE96 16'hC477
`define CUBE_LUT_BE95 16'hC475
`define CUBE_LUT_BE94 16'hC473
`define CUBE_LUT_BE93 16'hC471
`define CUBE_LUT_BE92 16'hC46F
`define CUBE_LUT_BE91 16'hC46D
`define CUBE_LUT_BE90 16'hC46A
`define CUBE_LUT_BE8F 16'hC468
`define CUBE_LUT_BE8E 16'hC466
`define CUBE_LUT_BE8D 16'hC464
`define CUBE_LUT_BE8C 16'hC462
`define CUBE_LUT_BE8B 16'hC460
`define CUBE_LUT_BE8A 16'hC45E
`define CUBE_LUT_BE89 16'hC45C
`define CUBE_LUT_BE88 16'hC45A
`define CUBE_LUT_BE87 16'hC458
`define CUBE_LUT_BE86 16'hC456
`define CUBE_LUT_BE85 16'hC454
`define CUBE_LUT_BE84 16'hC452
`define CUBE_LUT_BE83 16'hC450
`define CUBE_LUT_BE82 16'hC44E
`define CUBE_LUT_BE81 16'hC44C
`define CUBE_LUT_BE80 16'hC44A
`define CUBE_LUT_BE7F 16'hC449
`define CUBE_LUT_BE7E 16'hC447
`define CUBE_LUT_BE7D 16'hC445
`define CUBE_LUT_BE7C 16'hC443
`define CUBE_LUT_BE7B 16'hC441
`define CUBE_LUT_BE7A 16'hC43F
`define CUBE_LUT_BE79 16'hC43D
`define CUBE_LUT_BE78 16'hC43B
`define CUBE_LUT_BE77 16'hC439
`define CUBE_LUT_BE76 16'hC437
`define CUBE_LUT_BE75 16'hC435
`define CUBE_LUT_BE74 16'hC433
`define CUBE_LUT_BE73 16'hC431
`define CUBE_LUT_BE72 16'hC42F
`define CUBE_LUT_BE71 16'hC42D
`define CUBE_LUT_BE70 16'hC42B
`define CUBE_LUT_BE6F 16'hC429
`define CUBE_LUT_BE6E 16'hC427
`define CUBE_LUT_BE6D 16'hC425
`define CUBE_LUT_BE6C 16'hC423
`define CUBE_LUT_BE6B 16'hC421
`define CUBE_LUT_BE6A 16'hC420
`define CUBE_LUT_BE69 16'hC41E
`define CUBE_LUT_BE68 16'hC41C
`define CUBE_LUT_BE67 16'hC41A
`define CUBE_LUT_BE66 16'hC418
`define CUBE_LUT_BE65 16'hC416
`define CUBE_LUT_BE64 16'hC414
`define CUBE_LUT_BE63 16'hC412
`define CUBE_LUT_BE62 16'hC410
`define CUBE_LUT_BE61 16'hC40E
`define CUBE_LUT_BE60 16'hC40C
`define CUBE_LUT_BE5F 16'hC40A
`define CUBE_LUT_BE5E 16'hC409
`define CUBE_LUT_BE5D 16'hC407
`define CUBE_LUT_BE5C 16'hC405
`define CUBE_LUT_BE5B 16'hC403
`define CUBE_LUT_BE5A 16'hC401
`define CUBE_LUT_BE59 16'hC3FE
`define CUBE_LUT_BE58 16'hC3FA
`define CUBE_LUT_BE57 16'hC3F7
`define CUBE_LUT_BE56 16'hC3F3
`define CUBE_LUT_BE55 16'hC3EF
`define CUBE_LUT_BE54 16'hC3EB
`define CUBE_LUT_BE53 16'hC3E8
`define CUBE_LUT_BE52 16'hC3E4
`define CUBE_LUT_BE51 16'hC3E0
`define CUBE_LUT_BE50 16'hC3DC
`define CUBE_LUT_BE4F 16'hC3D9
`define CUBE_LUT_BE4E 16'hC3D5
`define CUBE_LUT_BE4D 16'hC3D1
`define CUBE_LUT_BE4C 16'hC3CD
`define CUBE_LUT_BE4B 16'hC3CA
`define CUBE_LUT_BE4A 16'hC3C6
`define CUBE_LUT_BE49 16'hC3C2
`define CUBE_LUT_BE48 16'hC3BF
`define CUBE_LUT_BE47 16'hC3BB
`define CUBE_LUT_BE46 16'hC3B7
`define CUBE_LUT_BE45 16'hC3B3
`define CUBE_LUT_BE44 16'hC3B0
`define CUBE_LUT_BE43 16'hC3AC
`define CUBE_LUT_BE42 16'hC3A8
`define CUBE_LUT_BE41 16'hC3A5
`define CUBE_LUT_BE40 16'hC3A1
`define CUBE_LUT_BE3F 16'hC39D
`define CUBE_LUT_BE3E 16'hC39A
`define CUBE_LUT_BE3D 16'hC396
`define CUBE_LUT_BE3C 16'hC393
`define CUBE_LUT_BE3B 16'hC38F
`define CUBE_LUT_BE3A 16'hC38B
`define CUBE_LUT_BE39 16'hC388
`define CUBE_LUT_BE38 16'hC384
`define CUBE_LUT_BE37 16'hC380
`define CUBE_LUT_BE36 16'hC37D
`define CUBE_LUT_BE35 16'hC379
`define CUBE_LUT_BE34 16'hC376
`define CUBE_LUT_BE33 16'hC372
`define CUBE_LUT_BE32 16'hC36E
`define CUBE_LUT_BE31 16'hC36B
`define CUBE_LUT_BE30 16'hC367
`define CUBE_LUT_BE2F 16'hC364
`define CUBE_LUT_BE2E 16'hC360
`define CUBE_LUT_BE2D 16'hC35C
`define CUBE_LUT_BE2C 16'hC359
`define CUBE_LUT_BE2B 16'hC355
`define CUBE_LUT_BE2A 16'hC352
`define CUBE_LUT_BE29 16'hC34E
`define CUBE_LUT_BE28 16'hC34B
`define CUBE_LUT_BE27 16'hC347
`define CUBE_LUT_BE26 16'hC343
`define CUBE_LUT_BE25 16'hC340
`define CUBE_LUT_BE24 16'hC33C
`define CUBE_LUT_BE23 16'hC339
`define CUBE_LUT_BE22 16'hC335
`define CUBE_LUT_BE21 16'hC332
`define CUBE_LUT_BE20 16'hC32E
`define CUBE_LUT_BE1F 16'hC32B
`define CUBE_LUT_BE1E 16'hC327
`define CUBE_LUT_BE1D 16'hC324
`define CUBE_LUT_BE1C 16'hC320
`define CUBE_LUT_BE1B 16'hC31D
`define CUBE_LUT_BE1A 16'hC319
`define CUBE_LUT_BE19 16'hC316
`define CUBE_LUT_BE18 16'hC312
`define CUBE_LUT_BE17 16'hC30F
`define CUBE_LUT_BE16 16'hC30B
`define CUBE_LUT_BE15 16'hC308
`define CUBE_LUT_BE14 16'hC304
`define CUBE_LUT_BE13 16'hC301
`define CUBE_LUT_BE12 16'hC2FD
`define CUBE_LUT_BE11 16'hC2FA
`define CUBE_LUT_BE10 16'hC2F7
`define CUBE_LUT_BE0F 16'hC2F3
`define CUBE_LUT_BE0E 16'hC2F0
`define CUBE_LUT_BE0D 16'hC2EC
`define CUBE_LUT_BE0C 16'hC2E9
`define CUBE_LUT_BE0B 16'hC2E5
`define CUBE_LUT_BE0A 16'hC2E2
`define CUBE_LUT_BE09 16'hC2DF
`define CUBE_LUT_BE08 16'hC2DB
`define CUBE_LUT_BE07 16'hC2D8
`define CUBE_LUT_BE06 16'hC2D4
`define CUBE_LUT_BE05 16'hC2D1
`define CUBE_LUT_BE04 16'hC2CE
`define CUBE_LUT_BE03 16'hC2CA
`define CUBE_LUT_BE02 16'hC2C7
`define CUBE_LUT_BE01 16'hC2C3
`define CUBE_LUT_BE00 16'hC2C0
`define CUBE_LUT_BDFF 16'hC2BD
`define CUBE_LUT_BDFE 16'hC2B9
`define CUBE_LUT_BDFD 16'hC2B6
`define CUBE_LUT_BDFC 16'hC2B3
`define CUBE_LUT_BDFB 16'hC2AF
`define CUBE_LUT_BDFA 16'hC2AC
`define CUBE_LUT_BDF9 16'hC2A8
`define CUBE_LUT_BDF8 16'hC2A5
`define CUBE_LUT_BDF7 16'hC2A2
`define CUBE_LUT_BDF6 16'hC29E
`define CUBE_LUT_BDF5 16'hC29B
`define CUBE_LUT_BDF4 16'hC298
`define CUBE_LUT_BDF3 16'hC294
`define CUBE_LUT_BDF2 16'hC291
`define CUBE_LUT_BDF1 16'hC28E
`define CUBE_LUT_BDF0 16'hC28B
`define CUBE_LUT_BDEF 16'hC287
`define CUBE_LUT_BDEE 16'hC284
`define CUBE_LUT_BDED 16'hC281
`define CUBE_LUT_BDEC 16'hC27D
`define CUBE_LUT_BDEB 16'hC27A
`define CUBE_LUT_BDEA 16'hC277
`define CUBE_LUT_BDE9 16'hC274
`define CUBE_LUT_BDE8 16'hC270
`define CUBE_LUT_BDE7 16'hC26D
`define CUBE_LUT_BDE6 16'hC26A
`define CUBE_LUT_BDE5 16'hC266
`define CUBE_LUT_BDE4 16'hC263
`define CUBE_LUT_BDE3 16'hC260
`define CUBE_LUT_BDE2 16'hC25D
`define CUBE_LUT_BDE1 16'hC259
`define CUBE_LUT_BDE0 16'hC256
`define CUBE_LUT_BDDF 16'hC253
`define CUBE_LUT_BDDE 16'hC250
`define CUBE_LUT_BDDD 16'hC24D
`define CUBE_LUT_BDDC 16'hC249
`define CUBE_LUT_BDDB 16'hC246
`define CUBE_LUT_BDDA 16'hC243
`define CUBE_LUT_BDD9 16'hC240
`define CUBE_LUT_BDD8 16'hC23C
`define CUBE_LUT_BDD7 16'hC239
`define CUBE_LUT_BDD6 16'hC236
`define CUBE_LUT_BDD5 16'hC233
`define CUBE_LUT_BDD4 16'hC230
`define CUBE_LUT_BDD3 16'hC22D
`define CUBE_LUT_BDD2 16'hC229
`define CUBE_LUT_BDD1 16'hC226
`define CUBE_LUT_BDD0 16'hC223
`define CUBE_LUT_BDCF 16'hC220
`define CUBE_LUT_BDCE 16'hC21D
`define CUBE_LUT_BDCD 16'hC21A
`define CUBE_LUT_BDCC 16'hC216
`define CUBE_LUT_BDCB 16'hC213
`define CUBE_LUT_BDCA 16'hC210
`define CUBE_LUT_BDC9 16'hC20D
`define CUBE_LUT_BDC8 16'hC20A
`define CUBE_LUT_BDC7 16'hC207
`define CUBE_LUT_BDC6 16'hC204
`define CUBE_LUT_BDC5 16'hC200
`define CUBE_LUT_BDC4 16'hC1FD
`define CUBE_LUT_BDC3 16'hC1FA
`define CUBE_LUT_BDC2 16'hC1F7
`define CUBE_LUT_BDC1 16'hC1F4
`define CUBE_LUT_BDC0 16'hC1F1
`define CUBE_LUT_BDBF 16'hC1EE
`define CUBE_LUT_BDBE 16'hC1EB
`define CUBE_LUT_BDBD 16'hC1E8
`define CUBE_LUT_BDBC 16'hC1E5
`define CUBE_LUT_BDBB 16'hC1E1
`define CUBE_LUT_BDBA 16'hC1DE
`define CUBE_LUT_BDB9 16'hC1DB
`define CUBE_LUT_BDB8 16'hC1D8
`define CUBE_LUT_BDB7 16'hC1D5
`define CUBE_LUT_BDB6 16'hC1D2
`define CUBE_LUT_BDB5 16'hC1CF
`define CUBE_LUT_BDB4 16'hC1CC
`define CUBE_LUT_BDB3 16'hC1C9
`define CUBE_LUT_BDB2 16'hC1C6
`define CUBE_LUT_BDB1 16'hC1C3
`define CUBE_LUT_BDB0 16'hC1C0
`define CUBE_LUT_BDAF 16'hC1BD
`define CUBE_LUT_BDAE 16'hC1BA
`define CUBE_LUT_BDAD 16'hC1B7
`define CUBE_LUT_BDAC 16'hC1B4
`define CUBE_LUT_BDAB 16'hC1B1
`define CUBE_LUT_BDAA 16'hC1AE
`define CUBE_LUT_BDA9 16'hC1AB
`define CUBE_LUT_BDA8 16'hC1A8
`define CUBE_LUT_BDA7 16'hC1A5
`define CUBE_LUT_BDA6 16'hC1A2
`define CUBE_LUT_BDA5 16'hC19F
`define CUBE_LUT_BDA4 16'hC19C
`define CUBE_LUT_BDA3 16'hC199
`define CUBE_LUT_BDA2 16'hC196
`define CUBE_LUT_BDA1 16'hC193
`define CUBE_LUT_BDA0 16'hC190
`define CUBE_LUT_BD9F 16'hC18D
`define CUBE_LUT_BD9E 16'hC18A
`define CUBE_LUT_BD9D 16'hC187
`define CUBE_LUT_BD9C 16'hC184
`define CUBE_LUT_BD9B 16'hC181
`define CUBE_LUT_BD9A 16'hC17E
`define CUBE_LUT_BD99 16'hC17B
`define CUBE_LUT_BD98 16'hC178
`define CUBE_LUT_BD97 16'hC175
`define CUBE_LUT_BD96 16'hC172
`define CUBE_LUT_BD95 16'hC16F
`define CUBE_LUT_BD94 16'hC16D
`define CUBE_LUT_BD93 16'hC16A
`define CUBE_LUT_BD92 16'hC167
`define CUBE_LUT_BD91 16'hC164
`define CUBE_LUT_BD90 16'hC161
`define CUBE_LUT_BD8F 16'hC15E
`define CUBE_LUT_BD8E 16'hC15B
`define CUBE_LUT_BD8D 16'hC158
`define CUBE_LUT_BD8C 16'hC155
`define CUBE_LUT_BD8B 16'hC152
`define CUBE_LUT_BD8A 16'hC150
`define CUBE_LUT_BD89 16'hC14D
`define CUBE_LUT_BD88 16'hC14A
`define CUBE_LUT_BD87 16'hC147
`define CUBE_LUT_BD86 16'hC144
`define CUBE_LUT_BD85 16'hC141
`define CUBE_LUT_BD84 16'hC13E
`define CUBE_LUT_BD83 16'hC13C
`define CUBE_LUT_BD82 16'hC139
`define CUBE_LUT_BD81 16'hC136
`define CUBE_LUT_BD80 16'hC133
`define CUBE_LUT_BD7F 16'hC130
`define CUBE_LUT_BD7E 16'hC12D
`define CUBE_LUT_BD7D 16'hC12B
`define CUBE_LUT_BD7C 16'hC128
`define CUBE_LUT_BD7B 16'hC125
`define CUBE_LUT_BD7A 16'hC122
`define CUBE_LUT_BD79 16'hC11F
`define CUBE_LUT_BD78 16'hC11C
`define CUBE_LUT_BD77 16'hC11A
`define CUBE_LUT_BD76 16'hC117
`define CUBE_LUT_BD75 16'hC114
`define CUBE_LUT_BD74 16'hC111
`define CUBE_LUT_BD73 16'hC10E
`define CUBE_LUT_BD72 16'hC10C
`define CUBE_LUT_BD71 16'hC109
`define CUBE_LUT_BD70 16'hC106
`define CUBE_LUT_BD6F 16'hC103
`define CUBE_LUT_BD6E 16'hC101
`define CUBE_LUT_BD6D 16'hC0FE
`define CUBE_LUT_BD6C 16'hC0FB
`define CUBE_LUT_BD6B 16'hC0F8
`define CUBE_LUT_BD6A 16'hC0F6
`define CUBE_LUT_BD69 16'hC0F3
`define CUBE_LUT_BD68 16'hC0F0
`define CUBE_LUT_BD67 16'hC0ED
`define CUBE_LUT_BD66 16'hC0EB
`define CUBE_LUT_BD65 16'hC0E8
`define CUBE_LUT_BD64 16'hC0E5
`define CUBE_LUT_BD63 16'hC0E2
`define CUBE_LUT_BD62 16'hC0E0
`define CUBE_LUT_BD61 16'hC0DD
`define CUBE_LUT_BD60 16'hC0DA
`define CUBE_LUT_BD5F 16'hC0D8
`define CUBE_LUT_BD5E 16'hC0D5
`define CUBE_LUT_BD5D 16'hC0D2
`define CUBE_LUT_BD5C 16'hC0CF
`define CUBE_LUT_BD5B 16'hC0CD
`define CUBE_LUT_BD5A 16'hC0CA
`define CUBE_LUT_BD59 16'hC0C7
`define CUBE_LUT_BD58 16'hC0C5
`define CUBE_LUT_BD57 16'hC0C2
`define CUBE_LUT_BD56 16'hC0BF
`define CUBE_LUT_BD55 16'hC0BD
`define CUBE_LUT_BD54 16'hC0BA
`define CUBE_LUT_BD53 16'hC0B7
`define CUBE_LUT_BD52 16'hC0B5
`define CUBE_LUT_BD51 16'hC0B2
`define CUBE_LUT_BD50 16'hC0AF
`define CUBE_LUT_BD4F 16'hC0AD
`define CUBE_LUT_BD4E 16'hC0AA
`define CUBE_LUT_BD4D 16'hC0A8
`define CUBE_LUT_BD4C 16'hC0A5
`define CUBE_LUT_BD4B 16'hC0A2
`define CUBE_LUT_BD4A 16'hC0A0
`define CUBE_LUT_BD49 16'hC09D
`define CUBE_LUT_BD48 16'hC09A
`define CUBE_LUT_BD47 16'hC098
`define CUBE_LUT_BD46 16'hC095
`define CUBE_LUT_BD45 16'hC093
`define CUBE_LUT_BD44 16'hC090
`define CUBE_LUT_BD43 16'hC08D
`define CUBE_LUT_BD42 16'hC08B
`define CUBE_LUT_BD41 16'hC088
`define CUBE_LUT_BD40 16'hC086
`define CUBE_LUT_BD3F 16'hC083
`define CUBE_LUT_BD3E 16'hC080
`define CUBE_LUT_BD3D 16'hC07E
`define CUBE_LUT_BD3C 16'hC07B
`define CUBE_LUT_BD3B 16'hC079
`define CUBE_LUT_BD3A 16'hC076
`define CUBE_LUT_BD39 16'hC074
`define CUBE_LUT_BD38 16'hC071
`define CUBE_LUT_BD37 16'hC06F
`define CUBE_LUT_BD36 16'hC06C
`define CUBE_LUT_BD35 16'hC069
`define CUBE_LUT_BD34 16'hC067
`define CUBE_LUT_BD33 16'hC064
`define CUBE_LUT_BD32 16'hC062
`define CUBE_LUT_BD31 16'hC05F
`define CUBE_LUT_BD30 16'hC05D
`define CUBE_LUT_BD2F 16'hC05A
`define CUBE_LUT_BD2E 16'hC058
`define CUBE_LUT_BD2D 16'hC055
`define CUBE_LUT_BD2C 16'hC053
`define CUBE_LUT_BD2B 16'hC050
`define CUBE_LUT_BD2A 16'hC04E
`define CUBE_LUT_BD29 16'hC04B
`define CUBE_LUT_BD28 16'hC049
`define CUBE_LUT_BD27 16'hC046
`define CUBE_LUT_BD26 16'hC044
`define CUBE_LUT_BD25 16'hC041
`define CUBE_LUT_BD24 16'hC03F
`define CUBE_LUT_BD23 16'hC03C
`define CUBE_LUT_BD22 16'hC03A
`define CUBE_LUT_BD21 16'hC037
`define CUBE_LUT_BD20 16'hC035
`define CUBE_LUT_BD1F 16'hC032
`define CUBE_LUT_BD1E 16'hC030
`define CUBE_LUT_BD1D 16'hC02E
`define CUBE_LUT_BD1C 16'hC02B
`define CUBE_LUT_BD1B 16'hC029
`define CUBE_LUT_BD1A 16'hC026
`define CUBE_LUT_BD19 16'hC024
`define CUBE_LUT_BD18 16'hC021
`define CUBE_LUT_BD17 16'hC01F
`define CUBE_LUT_BD16 16'hC01C
`define CUBE_LUT_BD15 16'hC01A
`define CUBE_LUT_BD14 16'hC018
`define CUBE_LUT_BD13 16'hC015
`define CUBE_LUT_BD12 16'hC013
`define CUBE_LUT_BD11 16'hC010
`define CUBE_LUT_BD10 16'hC00E
`define CUBE_LUT_BD0F 16'hC00C
`define CUBE_LUT_BD0E 16'hC009
`define CUBE_LUT_BD0D 16'hC007
`define CUBE_LUT_BD0C 16'hC004
`define CUBE_LUT_BD0B 16'hC002
`define CUBE_LUT_BD0A 16'hBFFF
`define CUBE_LUT_BD09 16'hBFFA
`define CUBE_LUT_BD08 16'hBFF6
`define CUBE_LUT_BD07 16'hBFF1
`define CUBE_LUT_BD06 16'hBFEC
`define CUBE_LUT_BD05 16'hBFE8
`define CUBE_LUT_BD04 16'hBFE3
`define CUBE_LUT_BD03 16'hBFDE
`define CUBE_LUT_BD02 16'hBFD9
`define CUBE_LUT_BD01 16'hBFD5
`define CUBE_LUT_BD00 16'hBFD0
`define CUBE_LUT_BCFF 16'hBFCB
`define CUBE_LUT_BCFE 16'hBFC7
`define CUBE_LUT_BCFD 16'hBFC2
`define CUBE_LUT_BCFC 16'hBFBD
`define CUBE_LUT_BCFB 16'hBFB9
`define CUBE_LUT_BCFA 16'hBFB4
`define CUBE_LUT_BCF9 16'hBFAF
`define CUBE_LUT_BCF8 16'hBFAB
`define CUBE_LUT_BCF7 16'hBFA6
`define CUBE_LUT_BCF6 16'hBFA1
`define CUBE_LUT_BCF5 16'hBF9D
`define CUBE_LUT_BCF4 16'hBF98
`define CUBE_LUT_BCF3 16'hBF94
`define CUBE_LUT_BCF2 16'hBF8F
`define CUBE_LUT_BCF1 16'hBF8B
`define CUBE_LUT_BCF0 16'hBF86
`define CUBE_LUT_BCEF 16'hBF81
`define CUBE_LUT_BCEE 16'hBF7D
`define CUBE_LUT_BCED 16'hBF78
`define CUBE_LUT_BCEC 16'hBF74
`define CUBE_LUT_BCEB 16'hBF6F
`define CUBE_LUT_BCEA 16'hBF6B
`define CUBE_LUT_BCE9 16'hBF66
`define CUBE_LUT_BCE8 16'hBF62
`define CUBE_LUT_BCE7 16'hBF5D
`define CUBE_LUT_BCE6 16'hBF59
`define CUBE_LUT_BCE5 16'hBF54
`define CUBE_LUT_BCE4 16'hBF50
`define CUBE_LUT_BCE3 16'hBF4B
`define CUBE_LUT_BCE2 16'hBF47
`define CUBE_LUT_BCE1 16'hBF42
`define CUBE_LUT_BCE0 16'hBF3E
`define CUBE_LUT_BCDF 16'hBF39
`define CUBE_LUT_BCDE 16'hBF35
`define CUBE_LUT_BCDD 16'hBF30
`define CUBE_LUT_BCDC 16'hBF2C
`define CUBE_LUT_BCDB 16'hBF28
`define CUBE_LUT_BCDA 16'hBF23
`define CUBE_LUT_BCD9 16'hBF1F
`define CUBE_LUT_BCD8 16'hBF1A
`define CUBE_LUT_BCD7 16'hBF16
`define CUBE_LUT_BCD6 16'hBF12
`define CUBE_LUT_BCD5 16'hBF0D
`define CUBE_LUT_BCD4 16'hBF09
`define CUBE_LUT_BCD3 16'hBF04
`define CUBE_LUT_BCD2 16'hBF00
`define CUBE_LUT_BCD1 16'hBEFC
`define CUBE_LUT_BCD0 16'hBEF7
`define CUBE_LUT_BCCF 16'hBEF3
`define CUBE_LUT_BCCE 16'hBEEF
`define CUBE_LUT_BCCD 16'hBEEA
`define CUBE_LUT_BCCC 16'hBEE6
`define CUBE_LUT_BCCB 16'hBEE2
`define CUBE_LUT_BCCA 16'hBEDD
`define CUBE_LUT_BCC9 16'hBED9
`define CUBE_LUT_BCC8 16'hBED5
`define CUBE_LUT_BCC7 16'hBED1
`define CUBE_LUT_BCC6 16'hBECC
`define CUBE_LUT_BCC5 16'hBEC8
`define CUBE_LUT_BCC4 16'hBEC4
`define CUBE_LUT_BCC3 16'hBEBF
`define CUBE_LUT_BCC2 16'hBEBB
`define CUBE_LUT_BCC1 16'hBEB7
`define CUBE_LUT_BCC0 16'hBEB3
`define CUBE_LUT_BCBF 16'hBEAF
`define CUBE_LUT_BCBE 16'hBEAA
`define CUBE_LUT_BCBD 16'hBEA6
`define CUBE_LUT_BCBC 16'hBEA2
`define CUBE_LUT_BCBB 16'hBE9E
`define CUBE_LUT_BCBA 16'hBE99
`define CUBE_LUT_BCB9 16'hBE95
`define CUBE_LUT_BCB8 16'hBE91
`define CUBE_LUT_BCB7 16'hBE8D
`define CUBE_LUT_BCB6 16'hBE89
`define CUBE_LUT_BCB5 16'hBE85
`define CUBE_LUT_BCB4 16'hBE80
`define CUBE_LUT_BCB3 16'hBE7C
`define CUBE_LUT_BCB2 16'hBE78
`define CUBE_LUT_BCB1 16'hBE74
`define CUBE_LUT_BCB0 16'hBE70
`define CUBE_LUT_BCAF 16'hBE6C
`define CUBE_LUT_BCAE 16'hBE68
`define CUBE_LUT_BCAD 16'hBE64
`define CUBE_LUT_BCAC 16'hBE60
`define CUBE_LUT_BCAB 16'hBE5B
`define CUBE_LUT_BCAA 16'hBE57
`define CUBE_LUT_BCA9 16'hBE53
`define CUBE_LUT_BCA8 16'hBE4F
`define CUBE_LUT_BCA7 16'hBE4B
`define CUBE_LUT_BCA6 16'hBE47
`define CUBE_LUT_BCA5 16'hBE43
`define CUBE_LUT_BCA4 16'hBE3F
`define CUBE_LUT_BCA3 16'hBE3B
`define CUBE_LUT_BCA2 16'hBE37
`define CUBE_LUT_BCA1 16'hBE33
`define CUBE_LUT_BCA0 16'hBE2F
`define CUBE_LUT_BC9F 16'hBE2B
`define CUBE_LUT_BC9E 16'hBE27
`define CUBE_LUT_BC9D 16'hBE23
`define CUBE_LUT_BC9C 16'hBE1F
`define CUBE_LUT_BC9B 16'hBE1B
`define CUBE_LUT_BC9A 16'hBE17
`define CUBE_LUT_BC99 16'hBE13
`define CUBE_LUT_BC98 16'hBE0F
`define CUBE_LUT_BC97 16'hBE0B
`define CUBE_LUT_BC96 16'hBE07
`define CUBE_LUT_BC95 16'hBE03
`define CUBE_LUT_BC94 16'hBDFF
`define CUBE_LUT_BC93 16'hBDFB
`define CUBE_LUT_BC92 16'hBDF7
`define CUBE_LUT_BC91 16'hBDF4
`define CUBE_LUT_BC90 16'hBDF0
`define CUBE_LUT_BC8F 16'hBDEC
`define CUBE_LUT_BC8E 16'hBDE8
`define CUBE_LUT_BC8D 16'hBDE4
`define CUBE_LUT_BC8C 16'hBDE0
`define CUBE_LUT_BC8B 16'hBDDC
`define CUBE_LUT_BC8A 16'hBDD8
`define CUBE_LUT_BC89 16'hBDD4
`define CUBE_LUT_BC88 16'hBDD1
`define CUBE_LUT_BC87 16'hBDCD
`define CUBE_LUT_BC86 16'hBDC9
`define CUBE_LUT_BC85 16'hBDC5
`define CUBE_LUT_BC84 16'hBDC1
`define CUBE_LUT_BC83 16'hBDBD
`define CUBE_LUT_BC82 16'hBDBA
`define CUBE_LUT_BC81 16'hBDB6
`define CUBE_LUT_BC80 16'hBDB2
`define CUBE_LUT_BC7F 16'hBDAE
`define CUBE_LUT_BC7E 16'hBDAA
`define CUBE_LUT_BC7D 16'hBDA7
`define CUBE_LUT_BC7C 16'hBDA3
`define CUBE_LUT_BC7B 16'hBD9F
`define CUBE_LUT_BC7A 16'hBD9B
`define CUBE_LUT_BC79 16'hBD98
`define CUBE_LUT_BC78 16'hBD94
`define CUBE_LUT_BC77 16'hBD90
`define CUBE_LUT_BC76 16'hBD8C
`define CUBE_LUT_BC75 16'hBD89
`define CUBE_LUT_BC74 16'hBD85
`define CUBE_LUT_BC73 16'hBD81
`define CUBE_LUT_BC72 16'hBD7D
`define CUBE_LUT_BC71 16'hBD7A
`define CUBE_LUT_BC70 16'hBD76
`define CUBE_LUT_BC6F 16'hBD72
`define CUBE_LUT_BC6E 16'hBD6F
`define CUBE_LUT_BC6D 16'hBD6B
`define CUBE_LUT_BC6C 16'hBD67
`define CUBE_LUT_BC6B 16'hBD64
`define CUBE_LUT_BC6A 16'hBD60
`define CUBE_LUT_BC69 16'hBD5C
`define CUBE_LUT_BC68 16'hBD59
`define CUBE_LUT_BC67 16'hBD55
`define CUBE_LUT_BC66 16'hBD51
`define CUBE_LUT_BC65 16'hBD4E
`define CUBE_LUT_BC64 16'hBD4A
`define CUBE_LUT_BC63 16'hBD47
`define CUBE_LUT_BC62 16'hBD43
`define CUBE_LUT_BC61 16'hBD3F
`define CUBE_LUT_BC60 16'hBD3C
`define CUBE_LUT_BC5F 16'hBD38
`define CUBE_LUT_BC5E 16'hBD35
`define CUBE_LUT_BC5D 16'hBD31
`define CUBE_LUT_BC5C 16'hBD2E
`define CUBE_LUT_BC5B 16'hBD2A
`define CUBE_LUT_BC5A 16'hBD26
`define CUBE_LUT_BC59 16'hBD23
`define CUBE_LUT_BC58 16'hBD1F
`define CUBE_LUT_BC57 16'hBD1C
`define CUBE_LUT_BC56 16'hBD18
`define CUBE_LUT_BC55 16'hBD15
`define CUBE_LUT_BC54 16'hBD11
`define CUBE_LUT_BC53 16'hBD0E
`define CUBE_LUT_BC52 16'hBD0A
`define CUBE_LUT_BC51 16'hBD07
`define CUBE_LUT_BC50 16'hBD03
`define CUBE_LUT_BC4F 16'hBD00
`define CUBE_LUT_BC4E 16'hBCFC
`define CUBE_LUT_BC4D 16'hBCF9
`define CUBE_LUT_BC4C 16'hBCF5
`define CUBE_LUT_BC4B 16'hBCF2
`define CUBE_LUT_BC4A 16'hBCEE
`define CUBE_LUT_BC49 16'hBCEB
`define CUBE_LUT_BC48 16'hBCE8
`define CUBE_LUT_BC47 16'hBCE4
`define CUBE_LUT_BC46 16'hBCE1
`define CUBE_LUT_BC45 16'hBCDD
`define CUBE_LUT_BC44 16'hBCDA
`define CUBE_LUT_BC43 16'hBCD6
`define CUBE_LUT_BC42 16'hBCD3
`define CUBE_LUT_BC41 16'hBCD0
`define CUBE_LUT_BC40 16'hBCCC
`define CUBE_LUT_BC3F 16'hBCC9
`define CUBE_LUT_BC3E 16'hBCC5
`define CUBE_LUT_BC3D 16'hBCC2
`define CUBE_LUT_BC3C 16'hBCBF
`define CUBE_LUT_BC3B 16'hBCBB
`define CUBE_LUT_BC3A 16'hBCB8
`define CUBE_LUT_BC39 16'hBCB5
`define CUBE_LUT_BC38 16'hBCB1
`define CUBE_LUT_BC37 16'hBCAE
`define CUBE_LUT_BC36 16'hBCAB
`define CUBE_LUT_BC35 16'hBCA7
`define CUBE_LUT_BC34 16'hBCA4
`define CUBE_LUT_BC33 16'hBCA1
`define CUBE_LUT_BC32 16'hBC9D
`define CUBE_LUT_BC31 16'hBC9A
`define CUBE_LUT_BC30 16'hBC97
`define CUBE_LUT_BC2F 16'hBC94
`define CUBE_LUT_BC2E 16'hBC90
`define CUBE_LUT_BC2D 16'hBC8D
`define CUBE_LUT_BC2C 16'hBC8A
`define CUBE_LUT_BC2B 16'hBC86
`define CUBE_LUT_BC2A 16'hBC83
`define CUBE_LUT_BC29 16'hBC80
`define CUBE_LUT_BC28 16'hBC7D
`define CUBE_LUT_BC27 16'hBC7A
`define CUBE_LUT_BC26 16'hBC76
`define CUBE_LUT_BC25 16'hBC73
`define CUBE_LUT_BC24 16'hBC70
`define CUBE_LUT_BC23 16'hBC6D
`define CUBE_LUT_BC22 16'hBC69
`define CUBE_LUT_BC21 16'hBC66
`define CUBE_LUT_BC20 16'hBC63
`define CUBE_LUT_BC1F 16'hBC60
`define CUBE_LUT_BC1E 16'hBC5D
`define CUBE_LUT_BC1D 16'hBC59
`define CUBE_LUT_BC1C 16'hBC56
`define CUBE_LUT_BC1B 16'hBC53
`define CUBE_LUT_BC1A 16'hBC50
`define CUBE_LUT_BC19 16'hBC4D
`define CUBE_LUT_BC18 16'hBC4A
`define CUBE_LUT_BC17 16'hBC47
`define CUBE_LUT_BC16 16'hBC43
`define CUBE_LUT_BC15 16'hBC40
`define CUBE_LUT_BC14 16'hBC3D
`define CUBE_LUT_BC13 16'hBC3A
`define CUBE_LUT_BC12 16'hBC37
`define CUBE_LUT_BC11 16'hBC34
`define CUBE_LUT_BC10 16'hBC31
`define CUBE_LUT_BC0F 16'hBC2E
`define CUBE_LUT_BC0E 16'hBC2B
`define CUBE_LUT_BC0D 16'hBC27
`define CUBE_LUT_BC0C 16'hBC24
`define CUBE_LUT_BC0B 16'hBC21
`define CUBE_LUT_BC0A 16'hBC1E
`define CUBE_LUT_BC09 16'hBC1B
`define CUBE_LUT_BC08 16'hBC18
`define CUBE_LUT_BC07 16'hBC15
`define CUBE_LUT_BC06 16'hBC12
`define CUBE_LUT_BC05 16'hBC0F
`define CUBE_LUT_BC04 16'hBC0C
`define CUBE_LUT_BC03 16'hBC09
`define CUBE_LUT_BC02 16'hBC06
`define CUBE_LUT_BC01 16'hBC03
`define CUBE_LUT_BC00 16'hBC00
`define CUBE_LUT_BBFF 16'hBBFD
`define CUBE_LUT_BBFE 16'hBBFA
`define CUBE_LUT_BBFD 16'hBBF7
`define CUBE_LUT_BBFC 16'hBBF4
`define CUBE_LUT_BBFB 16'hBBF1
`define CUBE_LUT_BBFA 16'hBBEE
`define CUBE_LUT_BBF9 16'hBBEB
`define CUBE_LUT_BBF8 16'hBBE8
`define CUBE_LUT_BBF7 16'hBBE5
`define CUBE_LUT_BBF6 16'hBBE2
`define CUBE_LUT_BBF5 16'hBBDF
`define CUBE_LUT_BBF4 16'hBBDC
`define CUBE_LUT_BBF3 16'hBBD9
`define CUBE_LUT_BBF2 16'hBBD6
`define CUBE_LUT_BBF1 16'hBBD3
`define CUBE_LUT_BBF0 16'hBBD0
`define CUBE_LUT_BBEF 16'hBBCD
`define CUBE_LUT_BBEE 16'hBBCA
`define CUBE_LUT_BBED 16'hBBC8
`define CUBE_LUT_BBEC 16'hBBC5
`define CUBE_LUT_BBEB 16'hBBC2
`define CUBE_LUT_BBEA 16'hBBBF
`define CUBE_LUT_BBE9 16'hBBBC
`define CUBE_LUT_BBE8 16'hBBB9
`define CUBE_LUT_BBE7 16'hBBB6
`define CUBE_LUT_BBE6 16'hBBB3
`define CUBE_LUT_BBE5 16'hBBB0
`define CUBE_LUT_BBE4 16'hBBAD
`define CUBE_LUT_BBE3 16'hBBAA
`define CUBE_LUT_BBE2 16'hBBA7
`define CUBE_LUT_BBE1 16'hBBA4
`define CUBE_LUT_BBE0 16'hBBA1
`define CUBE_LUT_BBDF 16'hBB9F
`define CUBE_LUT_BBDE 16'hBB9C
`define CUBE_LUT_BBDD 16'hBB99
`define CUBE_LUT_BBDC 16'hBB96
`define CUBE_LUT_BBDB 16'hBB93
`define CUBE_LUT_BBDA 16'hBB90
`define CUBE_LUT_BBD9 16'hBB8D
`define CUBE_LUT_BBD8 16'hBB8A
`define CUBE_LUT_BBD7 16'hBB87
`define CUBE_LUT_BBD6 16'hBB85
`define CUBE_LUT_BBD5 16'hBB82
`define CUBE_LUT_BBD4 16'hBB7F
`define CUBE_LUT_BBD3 16'hBB7C
`define CUBE_LUT_BBD2 16'hBB79
`define CUBE_LUT_BBD1 16'hBB76
`define CUBE_LUT_BBD0 16'hBB73
`define CUBE_LUT_BBCF 16'hBB70
`define CUBE_LUT_BBCE 16'hBB6E
`define CUBE_LUT_BBCD 16'hBB6B
`define CUBE_LUT_BBCC 16'hBB68
`define CUBE_LUT_BBCB 16'hBB65
`define CUBE_LUT_BBCA 16'hBB62
`define CUBE_LUT_BBC9 16'hBB5F
`define CUBE_LUT_BBC8 16'hBB5D
`define CUBE_LUT_BBC7 16'hBB5A
`define CUBE_LUT_BBC6 16'hBB57
`define CUBE_LUT_BBC5 16'hBB54
`define CUBE_LUT_BBC4 16'hBB51
`define CUBE_LUT_BBC3 16'hBB4E
`define CUBE_LUT_BBC2 16'hBB4C
`define CUBE_LUT_BBC1 16'hBB49
`define CUBE_LUT_BBC0 16'hBB46
`define CUBE_LUT_BBBF 16'hBB43
`define CUBE_LUT_BBBE 16'hBB40
`define CUBE_LUT_BBBD 16'hBB3E
`define CUBE_LUT_BBBC 16'hBB3B
`define CUBE_LUT_BBBB 16'hBB38
`define CUBE_LUT_BBBA 16'hBB35
`define CUBE_LUT_BBB9 16'hBB32
`define CUBE_LUT_BBB8 16'hBB30
`define CUBE_LUT_BBB7 16'hBB2D
`define CUBE_LUT_BBB6 16'hBB2A
`define CUBE_LUT_BBB5 16'hBB27
`define CUBE_LUT_BBB4 16'hBB24
`define CUBE_LUT_BBB3 16'hBB22
`define CUBE_LUT_BBB2 16'hBB1F
`define CUBE_LUT_BBB1 16'hBB1C
`define CUBE_LUT_BBB0 16'hBB19
`define CUBE_LUT_BBAF 16'hBB16
`define CUBE_LUT_BBAE 16'hBB14
`define CUBE_LUT_BBAD 16'hBB11
`define CUBE_LUT_BBAC 16'hBB0E
`define CUBE_LUT_BBAB 16'hBB0B
`define CUBE_LUT_BBAA 16'hBB09
`define CUBE_LUT_BBA9 16'hBB06
`define CUBE_LUT_BBA8 16'hBB03
`define CUBE_LUT_BBA7 16'hBB00
`define CUBE_LUT_BBA6 16'hBAFE
`define CUBE_LUT_BBA5 16'hBAFB
`define CUBE_LUT_BBA4 16'hBAF8
`define CUBE_LUT_BBA3 16'hBAF5
`define CUBE_LUT_BBA2 16'hBAF3
`define CUBE_LUT_BBA1 16'hBAF0
`define CUBE_LUT_BBA0 16'hBAED
`define CUBE_LUT_BB9F 16'hBAEB
`define CUBE_LUT_BB9E 16'hBAE8
`define CUBE_LUT_BB9D 16'hBAE5
`define CUBE_LUT_BB9C 16'hBAE2
`define CUBE_LUT_BB9B 16'hBAE0
`define CUBE_LUT_BB9A 16'hBADD
`define CUBE_LUT_BB99 16'hBADA
`define CUBE_LUT_BB98 16'hBAD8
`define CUBE_LUT_BB97 16'hBAD5
`define CUBE_LUT_BB96 16'hBAD2
`define CUBE_LUT_BB95 16'hBACF
`define CUBE_LUT_BB94 16'hBACD
`define CUBE_LUT_BB93 16'hBACA
`define CUBE_LUT_BB92 16'hBAC7
`define CUBE_LUT_BB91 16'hBAC5
`define CUBE_LUT_BB90 16'hBAC2
`define CUBE_LUT_BB8F 16'hBABF
`define CUBE_LUT_BB8E 16'hBABD
`define CUBE_LUT_BB8D 16'hBABA
`define CUBE_LUT_BB8C 16'hBAB7
`define CUBE_LUT_BB8B 16'hBAB5
`define CUBE_LUT_BB8A 16'hBAB2
`define CUBE_LUT_BB89 16'hBAAF
`define CUBE_LUT_BB88 16'hBAAD
`define CUBE_LUT_BB87 16'hBAAA
`define CUBE_LUT_BB86 16'hBAA7
`define CUBE_LUT_BB85 16'hBAA5
`define CUBE_LUT_BB84 16'hBAA2
`define CUBE_LUT_BB83 16'hBA9F
`define CUBE_LUT_BB82 16'hBA9D
`define CUBE_LUT_BB81 16'hBA9A
`define CUBE_LUT_BB80 16'hBA98
`define CUBE_LUT_BB7F 16'hBA95
`define CUBE_LUT_BB7E 16'hBA92
`define CUBE_LUT_BB7D 16'hBA90
`define CUBE_LUT_BB7C 16'hBA8D
`define CUBE_LUT_BB7B 16'hBA8A
`define CUBE_LUT_BB7A 16'hBA88
`define CUBE_LUT_BB79 16'hBA85
`define CUBE_LUT_BB78 16'hBA82
`define CUBE_LUT_BB77 16'hBA80
`define CUBE_LUT_BB76 16'hBA7D
`define CUBE_LUT_BB75 16'hBA7B
`define CUBE_LUT_BB74 16'hBA78
`define CUBE_LUT_BB73 16'hBA75
`define CUBE_LUT_BB72 16'hBA73
`define CUBE_LUT_BB71 16'hBA70
`define CUBE_LUT_BB70 16'hBA6E
`define CUBE_LUT_BB6F 16'hBA6B
`define CUBE_LUT_BB6E 16'hBA68
`define CUBE_LUT_BB6D 16'hBA66
`define CUBE_LUT_BB6C 16'hBA63
`define CUBE_LUT_BB6B 16'hBA61
`define CUBE_LUT_BB6A 16'hBA5E
`define CUBE_LUT_BB69 16'hBA5C
`define CUBE_LUT_BB68 16'hBA59
`define CUBE_LUT_BB67 16'hBA56
`define CUBE_LUT_BB66 16'hBA54
`define CUBE_LUT_BB65 16'hBA51
`define CUBE_LUT_BB64 16'hBA4F
`define CUBE_LUT_BB63 16'hBA4C
`define CUBE_LUT_BB62 16'hBA4A
`define CUBE_LUT_BB61 16'hBA47
`define CUBE_LUT_BB60 16'hBA45
`define CUBE_LUT_BB5F 16'hBA42
`define CUBE_LUT_BB5E 16'hBA3F
`define CUBE_LUT_BB5D 16'hBA3D
`define CUBE_LUT_BB5C 16'hBA3A
`define CUBE_LUT_BB5B 16'hBA38
`define CUBE_LUT_BB5A 16'hBA35
`define CUBE_LUT_BB59 16'hBA33
`define CUBE_LUT_BB58 16'hBA30
`define CUBE_LUT_BB57 16'hBA2E
`define CUBE_LUT_BB56 16'hBA2B
`define CUBE_LUT_BB55 16'hBA29
`define CUBE_LUT_BB54 16'hBA26
`define CUBE_LUT_BB53 16'hBA24
`define CUBE_LUT_BB52 16'hBA21
`define CUBE_LUT_BB51 16'hBA1F
`define CUBE_LUT_BB50 16'hBA1C
`define CUBE_LUT_BB4F 16'hBA1A
`define CUBE_LUT_BB4E 16'hBA17
`define CUBE_LUT_BB4D 16'hBA15
`define CUBE_LUT_BB4C 16'hBA12
`define CUBE_LUT_BB4B 16'hBA10
`define CUBE_LUT_BB4A 16'hBA0D
`define CUBE_LUT_BB49 16'hBA0B
`define CUBE_LUT_BB48 16'hBA08
`define CUBE_LUT_BB47 16'hBA06
`define CUBE_LUT_BB46 16'hBA03
`define CUBE_LUT_BB45 16'hBA01
`define CUBE_LUT_BB44 16'hB9FE
`define CUBE_LUT_BB43 16'hB9FC
`define CUBE_LUT_BB42 16'hB9F9
`define CUBE_LUT_BB41 16'hB9F7
`define CUBE_LUT_BB40 16'hB9F4
`define CUBE_LUT_BB3F 16'hB9F2
`define CUBE_LUT_BB3E 16'hB9EF
`define CUBE_LUT_BB3D 16'hB9ED
`define CUBE_LUT_BB3C 16'hB9EA
`define CUBE_LUT_BB3B 16'hB9E8
`define CUBE_LUT_BB3A 16'hB9E6
`define CUBE_LUT_BB39 16'hB9E3
`define CUBE_LUT_BB38 16'hB9E1
`define CUBE_LUT_BB37 16'hB9DE
`define CUBE_LUT_BB36 16'hB9DC
`define CUBE_LUT_BB35 16'hB9D9
`define CUBE_LUT_BB34 16'hB9D7
`define CUBE_LUT_BB33 16'hB9D5
`define CUBE_LUT_BB32 16'hB9D2
`define CUBE_LUT_BB31 16'hB9D0
`define CUBE_LUT_BB30 16'hB9CD
`define CUBE_LUT_BB2F 16'hB9CB
`define CUBE_LUT_BB2E 16'hB9C8
`define CUBE_LUT_BB2D 16'hB9C6
`define CUBE_LUT_BB2C 16'hB9C4
`define CUBE_LUT_BB2B 16'hB9C1
`define CUBE_LUT_BB2A 16'hB9BF
`define CUBE_LUT_BB29 16'hB9BC
`define CUBE_LUT_BB28 16'hB9BA
`define CUBE_LUT_BB27 16'hB9B8
`define CUBE_LUT_BB26 16'hB9B5
`define CUBE_LUT_BB25 16'hB9B3
`define CUBE_LUT_BB24 16'hB9B0
`define CUBE_LUT_BB23 16'hB9AE
`define CUBE_LUT_BB22 16'hB9AC
`define CUBE_LUT_BB21 16'hB9A9
`define CUBE_LUT_BB20 16'hB9A7
`define CUBE_LUT_BB1F 16'hB9A4
`define CUBE_LUT_BB1E 16'hB9A2
`define CUBE_LUT_BB1D 16'hB9A0
`define CUBE_LUT_BB1C 16'hB99D
`define CUBE_LUT_BB1B 16'hB99B
`define CUBE_LUT_BB1A 16'hB999
`define CUBE_LUT_BB19 16'hB996
`define CUBE_LUT_BB18 16'hB994
`define CUBE_LUT_BB17 16'hB992
`define CUBE_LUT_BB16 16'hB98F
`define CUBE_LUT_BB15 16'hB98D
`define CUBE_LUT_BB14 16'hB98A
`define CUBE_LUT_BB13 16'hB988
`define CUBE_LUT_BB12 16'hB986
`define CUBE_LUT_BB11 16'hB983
`define CUBE_LUT_BB10 16'hB981
`define CUBE_LUT_BB0F 16'hB97F
`define CUBE_LUT_BB0E 16'hB97C
`define CUBE_LUT_BB0D 16'hB97A
`define CUBE_LUT_BB0C 16'hB978
`define CUBE_LUT_BB0B 16'hB975
`define CUBE_LUT_BB0A 16'hB973
`define CUBE_LUT_BB09 16'hB971
`define CUBE_LUT_BB08 16'hB96E
`define CUBE_LUT_BB07 16'hB96C
`define CUBE_LUT_BB06 16'hB96A
`define CUBE_LUT_BB05 16'hB968
`define CUBE_LUT_BB04 16'hB965
`define CUBE_LUT_BB03 16'hB963
`define CUBE_LUT_BB02 16'hB961
`define CUBE_LUT_BB01 16'hB95E
`define CUBE_LUT_BB00 16'hB95C
`define CUBE_LUT_BAFF 16'hB95A
`define CUBE_LUT_BAFE 16'hB957
`define CUBE_LUT_BAFD 16'hB955
`define CUBE_LUT_BAFC 16'hB953
`define CUBE_LUT_BAFB 16'hB951
`define CUBE_LUT_BAFA 16'hB94E
`define CUBE_LUT_BAF9 16'hB94C
`define CUBE_LUT_BAF8 16'hB94A
`define CUBE_LUT_BAF7 16'hB947
`define CUBE_LUT_BAF6 16'hB945
`define CUBE_LUT_BAF5 16'hB943
`define CUBE_LUT_BAF4 16'hB941
`define CUBE_LUT_BAF3 16'hB93E
`define CUBE_LUT_BAF2 16'hB93C
`define CUBE_LUT_BAF1 16'hB93A
`define CUBE_LUT_BAF0 16'hB938
`define CUBE_LUT_BAEF 16'hB935
`define CUBE_LUT_BAEE 16'hB933
`define CUBE_LUT_BAED 16'hB931
`define CUBE_LUT_BAEC 16'hB92F
`define CUBE_LUT_BAEB 16'hB92C
`define CUBE_LUT_BAEA 16'hB92A
`define CUBE_LUT_BAE9 16'hB928
`define CUBE_LUT_BAE8 16'hB926
`define CUBE_LUT_BAE7 16'hB923
`define CUBE_LUT_BAE6 16'hB921
`define CUBE_LUT_BAE5 16'hB91F
`define CUBE_LUT_BAE4 16'hB91D
`define CUBE_LUT_BAE3 16'hB91A
`define CUBE_LUT_BAE2 16'hB918
`define CUBE_LUT_BAE1 16'hB916
`define CUBE_LUT_BAE0 16'hB914
`define CUBE_LUT_BADF 16'hB912
`define CUBE_LUT_BADE 16'hB90F
`define CUBE_LUT_BADD 16'hB90D
`define CUBE_LUT_BADC 16'hB90B
`define CUBE_LUT_BADB 16'hB909
`define CUBE_LUT_BADA 16'hB907
`define CUBE_LUT_BAD9 16'hB904
`define CUBE_LUT_BAD8 16'hB902
`define CUBE_LUT_BAD7 16'hB900
`define CUBE_LUT_BAD6 16'hB8FE
`define CUBE_LUT_BAD5 16'hB8FC
`define CUBE_LUT_BAD4 16'hB8F9
`define CUBE_LUT_BAD3 16'hB8F7
`define CUBE_LUT_BAD2 16'hB8F5
`define CUBE_LUT_BAD1 16'hB8F3
`define CUBE_LUT_BAD0 16'hB8F1
`define CUBE_LUT_BACF 16'hB8EF
`define CUBE_LUT_BACE 16'hB8EC
`define CUBE_LUT_BACD 16'hB8EA
`define CUBE_LUT_BACC 16'hB8E8
`define CUBE_LUT_BACB 16'hB8E6
`define CUBE_LUT_BACA 16'hB8E4
`define CUBE_LUT_BAC9 16'hB8E2
`define CUBE_LUT_BAC8 16'hB8DF
`define CUBE_LUT_BAC7 16'hB8DD
`define CUBE_LUT_BAC6 16'hB8DB
`define CUBE_LUT_BAC5 16'hB8D9
`define CUBE_LUT_BAC4 16'hB8D7
`define CUBE_LUT_BAC3 16'hB8D5
`define CUBE_LUT_BAC2 16'hB8D2
`define CUBE_LUT_BAC1 16'hB8D0
`define CUBE_LUT_BAC0 16'hB8CE
`define CUBE_LUT_BABF 16'hB8CC
`define CUBE_LUT_BABE 16'hB8CA
`define CUBE_LUT_BABD 16'hB8C8
`define CUBE_LUT_BABC 16'hB8C6
`define CUBE_LUT_BABB 16'hB8C4
`define CUBE_LUT_BABA 16'hB8C1
`define CUBE_LUT_BAB9 16'hB8BF
`define CUBE_LUT_BAB8 16'hB8BD
`define CUBE_LUT_BAB7 16'hB8BB
`define CUBE_LUT_BAB6 16'hB8B9
`define CUBE_LUT_BAB5 16'hB8B7
`define CUBE_LUT_BAB4 16'hB8B5
`define CUBE_LUT_BAB3 16'hB8B3
`define CUBE_LUT_BAB2 16'hB8B1
`define CUBE_LUT_BAB1 16'hB8AE
`define CUBE_LUT_BAB0 16'hB8AC
`define CUBE_LUT_BAAF 16'hB8AA
`define CUBE_LUT_BAAE 16'hB8A8
`define CUBE_LUT_BAAD 16'hB8A6
`define CUBE_LUT_BAAC 16'hB8A4
`define CUBE_LUT_BAAB 16'hB8A2
`define CUBE_LUT_BAAA 16'hB8A0
`define CUBE_LUT_BAA9 16'hB89E
`define CUBE_LUT_BAA8 16'hB89C
`define CUBE_LUT_BAA7 16'hB89A
`define CUBE_LUT_BAA6 16'hB897
`define CUBE_LUT_BAA5 16'hB895
`define CUBE_LUT_BAA4 16'hB893
`define CUBE_LUT_BAA3 16'hB891
`define CUBE_LUT_BAA2 16'hB88F
`define CUBE_LUT_BAA1 16'hB88D
`define CUBE_LUT_BAA0 16'hB88B
`define CUBE_LUT_BA9F 16'hB889
`define CUBE_LUT_BA9E 16'hB887
`define CUBE_LUT_BA9D 16'hB885
`define CUBE_LUT_BA9C 16'hB883
`define CUBE_LUT_BA9B 16'hB881
`define CUBE_LUT_BA9A 16'hB87F
`define CUBE_LUT_BA99 16'hB87D
`define CUBE_LUT_BA98 16'hB87B
`define CUBE_LUT_BA97 16'hB879
`define CUBE_LUT_BA96 16'hB877
`define CUBE_LUT_BA95 16'hB875
`define CUBE_LUT_BA94 16'hB873
`define CUBE_LUT_BA93 16'hB871
`define CUBE_LUT_BA92 16'hB86F
`define CUBE_LUT_BA91 16'hB86D
`define CUBE_LUT_BA90 16'hB86A
`define CUBE_LUT_BA8F 16'hB868
`define CUBE_LUT_BA8E 16'hB866
`define CUBE_LUT_BA8D 16'hB864
`define CUBE_LUT_BA8C 16'hB862
`define CUBE_LUT_BA8B 16'hB860
`define CUBE_LUT_BA8A 16'hB85E
`define CUBE_LUT_BA89 16'hB85C
`define CUBE_LUT_BA88 16'hB85A
`define CUBE_LUT_BA87 16'hB858
`define CUBE_LUT_BA86 16'hB856
`define CUBE_LUT_BA85 16'hB854
`define CUBE_LUT_BA84 16'hB852
`define CUBE_LUT_BA83 16'hB850
`define CUBE_LUT_BA82 16'hB84E
`define CUBE_LUT_BA81 16'hB84C
`define CUBE_LUT_BA80 16'hB84A
`define CUBE_LUT_BA7F 16'hB849
`define CUBE_LUT_BA7E 16'hB847
`define CUBE_LUT_BA7D 16'hB845
`define CUBE_LUT_BA7C 16'hB843
`define CUBE_LUT_BA7B 16'hB841
`define CUBE_LUT_BA7A 16'hB83F
`define CUBE_LUT_BA79 16'hB83D
`define CUBE_LUT_BA78 16'hB83B
`define CUBE_LUT_BA77 16'hB839
`define CUBE_LUT_BA76 16'hB837
`define CUBE_LUT_BA75 16'hB835
`define CUBE_LUT_BA74 16'hB833
`define CUBE_LUT_BA73 16'hB831
`define CUBE_LUT_BA72 16'hB82F
`define CUBE_LUT_BA71 16'hB82D
`define CUBE_LUT_BA70 16'hB82B
`define CUBE_LUT_BA6F 16'hB829
`define CUBE_LUT_BA6E 16'hB827
`define CUBE_LUT_BA6D 16'hB825
`define CUBE_LUT_BA6C 16'hB823
`define CUBE_LUT_BA6B 16'hB821
`define CUBE_LUT_BA6A 16'hB820
`define CUBE_LUT_BA69 16'hB81E
`define CUBE_LUT_BA68 16'hB81C
`define CUBE_LUT_BA67 16'hB81A
`define CUBE_LUT_BA66 16'hB818
`define CUBE_LUT_BA65 16'hB816
`define CUBE_LUT_BA64 16'hB814
`define CUBE_LUT_BA63 16'hB812
`define CUBE_LUT_BA62 16'hB810
`define CUBE_LUT_BA61 16'hB80E
`define CUBE_LUT_BA60 16'hB80C
`define CUBE_LUT_BA5F 16'hB80A
`define CUBE_LUT_BA5E 16'hB809
`define CUBE_LUT_BA5D 16'hB807
`define CUBE_LUT_BA5C 16'hB805
`define CUBE_LUT_BA5B 16'hB803
`define CUBE_LUT_BA5A 16'hB801
`define CUBE_LUT_BA59 16'hB7FE
`define CUBE_LUT_BA58 16'hB7FA
`define CUBE_LUT_BA57 16'hB7F7
`define CUBE_LUT_BA56 16'hB7F3
`define CUBE_LUT_BA55 16'hB7EF
`define CUBE_LUT_BA54 16'hB7EB
`define CUBE_LUT_BA53 16'hB7E8
`define CUBE_LUT_BA52 16'hB7E4
`define CUBE_LUT_BA51 16'hB7E0
`define CUBE_LUT_BA50 16'hB7DC
`define CUBE_LUT_BA4F 16'hB7D9
`define CUBE_LUT_BA4E 16'hB7D5
`define CUBE_LUT_BA4D 16'hB7D1
`define CUBE_LUT_BA4C 16'hB7CD
`define CUBE_LUT_BA4B 16'hB7CA
`define CUBE_LUT_BA4A 16'hB7C6
`define CUBE_LUT_BA49 16'hB7C2
`define CUBE_LUT_BA48 16'hB7BF
`define CUBE_LUT_BA47 16'hB7BB
`define CUBE_LUT_BA46 16'hB7B7
`define CUBE_LUT_BA45 16'hB7B3
`define CUBE_LUT_BA44 16'hB7B0
`define CUBE_LUT_BA43 16'hB7AC
`define CUBE_LUT_BA42 16'hB7A8
`define CUBE_LUT_BA41 16'hB7A5
`define CUBE_LUT_BA40 16'hB7A1
`define CUBE_LUT_BA3F 16'hB79D
`define CUBE_LUT_BA3E 16'hB79A
`define CUBE_LUT_BA3D 16'hB796
`define CUBE_LUT_BA3C 16'hB793
`define CUBE_LUT_BA3B 16'hB78F
`define CUBE_LUT_BA3A 16'hB78B
`define CUBE_LUT_BA39 16'hB788
`define CUBE_LUT_BA38 16'hB784
`define CUBE_LUT_BA37 16'hB780
`define CUBE_LUT_BA36 16'hB77D
`define CUBE_LUT_BA35 16'hB779
`define CUBE_LUT_BA34 16'hB776
`define CUBE_LUT_BA33 16'hB772
`define CUBE_LUT_BA32 16'hB76E
`define CUBE_LUT_BA31 16'hB76B
`define CUBE_LUT_BA30 16'hB767
`define CUBE_LUT_BA2F 16'hB764
`define CUBE_LUT_BA2E 16'hB760
`define CUBE_LUT_BA2D 16'hB75C
`define CUBE_LUT_BA2C 16'hB759
`define CUBE_LUT_BA2B 16'hB755
`define CUBE_LUT_BA2A 16'hB752
`define CUBE_LUT_BA29 16'hB74E
`define CUBE_LUT_BA28 16'hB74B
`define CUBE_LUT_BA27 16'hB747
`define CUBE_LUT_BA26 16'hB743
`define CUBE_LUT_BA25 16'hB740
`define CUBE_LUT_BA24 16'hB73C
`define CUBE_LUT_BA23 16'hB739
`define CUBE_LUT_BA22 16'hB735
`define CUBE_LUT_BA21 16'hB732
`define CUBE_LUT_BA20 16'hB72E
`define CUBE_LUT_BA1F 16'hB72B
`define CUBE_LUT_BA1E 16'hB727
`define CUBE_LUT_BA1D 16'hB724
`define CUBE_LUT_BA1C 16'hB720
`define CUBE_LUT_BA1B 16'hB71D
`define CUBE_LUT_BA1A 16'hB719
`define CUBE_LUT_BA19 16'hB716
`define CUBE_LUT_BA18 16'hB712
`define CUBE_LUT_BA17 16'hB70F
`define CUBE_LUT_BA16 16'hB70B
`define CUBE_LUT_BA15 16'hB708
`define CUBE_LUT_BA14 16'hB704
`define CUBE_LUT_BA13 16'hB701
`define CUBE_LUT_BA12 16'hB6FD
`define CUBE_LUT_BA11 16'hB6FA
`define CUBE_LUT_BA10 16'hB6F7
`define CUBE_LUT_BA0F 16'hB6F3
`define CUBE_LUT_BA0E 16'hB6F0
`define CUBE_LUT_BA0D 16'hB6EC
`define CUBE_LUT_BA0C 16'hB6E9
`define CUBE_LUT_BA0B 16'hB6E5
`define CUBE_LUT_BA0A 16'hB6E2
`define CUBE_LUT_BA09 16'hB6DF
`define CUBE_LUT_BA08 16'hB6DB
`define CUBE_LUT_BA07 16'hB6D8
`define CUBE_LUT_BA06 16'hB6D4
`define CUBE_LUT_BA05 16'hB6D1
`define CUBE_LUT_BA04 16'hB6CE
`define CUBE_LUT_BA03 16'hB6CA
`define CUBE_LUT_BA02 16'hB6C7
`define CUBE_LUT_BA01 16'hB6C3
`define CUBE_LUT_BA00 16'hB6C0
`define CUBE_LUT_B9FF 16'hB6BD
`define CUBE_LUT_B9FE 16'hB6B9
`define CUBE_LUT_B9FD 16'hB6B6
`define CUBE_LUT_B9FC 16'hB6B3
`define CUBE_LUT_B9FB 16'hB6AF
`define CUBE_LUT_B9FA 16'hB6AC
`define CUBE_LUT_B9F9 16'hB6A8
`define CUBE_LUT_B9F8 16'hB6A5
`define CUBE_LUT_B9F7 16'hB6A2
`define CUBE_LUT_B9F6 16'hB69E
`define CUBE_LUT_B9F5 16'hB69B
`define CUBE_LUT_B9F4 16'hB698
`define CUBE_LUT_B9F3 16'hB694
`define CUBE_LUT_B9F2 16'hB691
`define CUBE_LUT_B9F1 16'hB68E
`define CUBE_LUT_B9F0 16'hB68B
`define CUBE_LUT_B9EF 16'hB687
`define CUBE_LUT_B9EE 16'hB684
`define CUBE_LUT_B9ED 16'hB681
`define CUBE_LUT_B9EC 16'hB67D
`define CUBE_LUT_B9EB 16'hB67A
`define CUBE_LUT_B9EA 16'hB677
`define CUBE_LUT_B9E9 16'hB674
`define CUBE_LUT_B9E8 16'hB670
`define CUBE_LUT_B9E7 16'hB66D
`define CUBE_LUT_B9E6 16'hB66A
`define CUBE_LUT_B9E5 16'hB666
`define CUBE_LUT_B9E4 16'hB663
`define CUBE_LUT_B9E3 16'hB660
`define CUBE_LUT_B9E2 16'hB65D
`define CUBE_LUT_B9E1 16'hB659
`define CUBE_LUT_B9E0 16'hB656
`define CUBE_LUT_B9DF 16'hB653
`define CUBE_LUT_B9DE 16'hB650
`define CUBE_LUT_B9DD 16'hB64D
`define CUBE_LUT_B9DC 16'hB649
`define CUBE_LUT_B9DB 16'hB646
`define CUBE_LUT_B9DA 16'hB643
`define CUBE_LUT_B9D9 16'hB640
`define CUBE_LUT_B9D8 16'hB63C
`define CUBE_LUT_B9D7 16'hB639
`define CUBE_LUT_B9D6 16'hB636
`define CUBE_LUT_B9D5 16'hB633
`define CUBE_LUT_B9D4 16'hB630
`define CUBE_LUT_B9D3 16'hB62D
`define CUBE_LUT_B9D2 16'hB629
`define CUBE_LUT_B9D1 16'hB626
`define CUBE_LUT_B9D0 16'hB623
`define CUBE_LUT_B9CF 16'hB620
`define CUBE_LUT_B9CE 16'hB61D
`define CUBE_LUT_B9CD 16'hB61A
`define CUBE_LUT_B9CC 16'hB616
`define CUBE_LUT_B9CB 16'hB613
`define CUBE_LUT_B9CA 16'hB610
`define CUBE_LUT_B9C9 16'hB60D
`define CUBE_LUT_B9C8 16'hB60A
`define CUBE_LUT_B9C7 16'hB607
`define CUBE_LUT_B9C6 16'hB604
`define CUBE_LUT_B9C5 16'hB600
`define CUBE_LUT_B9C4 16'hB5FD
`define CUBE_LUT_B9C3 16'hB5FA
`define CUBE_LUT_B9C2 16'hB5F7
`define CUBE_LUT_B9C1 16'hB5F4
`define CUBE_LUT_B9C0 16'hB5F1
`define CUBE_LUT_B9BF 16'hB5EE
`define CUBE_LUT_B9BE 16'hB5EB
`define CUBE_LUT_B9BD 16'hB5E8
`define CUBE_LUT_B9BC 16'hB5E5
`define CUBE_LUT_B9BB 16'hB5E1
`define CUBE_LUT_B9BA 16'hB5DE
`define CUBE_LUT_B9B9 16'hB5DB
`define CUBE_LUT_B9B8 16'hB5D8
`define CUBE_LUT_B9B7 16'hB5D5
`define CUBE_LUT_B9B6 16'hB5D2
`define CUBE_LUT_B9B5 16'hB5CF
`define CUBE_LUT_B9B4 16'hB5CC
`define CUBE_LUT_B9B3 16'hB5C9
`define CUBE_LUT_B9B2 16'hB5C6
`define CUBE_LUT_B9B1 16'hB5C3
`define CUBE_LUT_B9B0 16'hB5C0
`define CUBE_LUT_B9AF 16'hB5BD
`define CUBE_LUT_B9AE 16'hB5BA
`define CUBE_LUT_B9AD 16'hB5B7
`define CUBE_LUT_B9AC 16'hB5B4
`define CUBE_LUT_B9AB 16'hB5B1
`define CUBE_LUT_B9AA 16'hB5AE
`define CUBE_LUT_B9A9 16'hB5AB
`define CUBE_LUT_B9A8 16'hB5A8
`define CUBE_LUT_B9A7 16'hB5A5
`define CUBE_LUT_B9A6 16'hB5A2
`define CUBE_LUT_B9A5 16'hB59F
`define CUBE_LUT_B9A4 16'hB59C
`define CUBE_LUT_B9A3 16'hB599
`define CUBE_LUT_B9A2 16'hB596
`define CUBE_LUT_B9A1 16'hB593
`define CUBE_LUT_B9A0 16'hB590
`define CUBE_LUT_B99F 16'hB58D
`define CUBE_LUT_B99E 16'hB58A
`define CUBE_LUT_B99D 16'hB587
`define CUBE_LUT_B99C 16'hB584
`define CUBE_LUT_B99B 16'hB581
`define CUBE_LUT_B99A 16'hB57E
`define CUBE_LUT_B999 16'hB57B
`define CUBE_LUT_B998 16'hB578
`define CUBE_LUT_B997 16'hB575
`define CUBE_LUT_B996 16'hB572
`define CUBE_LUT_B995 16'hB56F
`define CUBE_LUT_B994 16'hB56D
`define CUBE_LUT_B993 16'hB56A
`define CUBE_LUT_B992 16'hB567
`define CUBE_LUT_B991 16'hB564
`define CUBE_LUT_B990 16'hB561
`define CUBE_LUT_B98F 16'hB55E
`define CUBE_LUT_B98E 16'hB55B
`define CUBE_LUT_B98D 16'hB558
`define CUBE_LUT_B98C 16'hB555
`define CUBE_LUT_B98B 16'hB552
`define CUBE_LUT_B98A 16'hB550
`define CUBE_LUT_B989 16'hB54D
`define CUBE_LUT_B988 16'hB54A
`define CUBE_LUT_B987 16'hB547
`define CUBE_LUT_B986 16'hB544
`define CUBE_LUT_B985 16'hB541
`define CUBE_LUT_B984 16'hB53E
`define CUBE_LUT_B983 16'hB53C
`define CUBE_LUT_B982 16'hB539
`define CUBE_LUT_B981 16'hB536
`define CUBE_LUT_B980 16'hB533
`define CUBE_LUT_B97F 16'hB530
`define CUBE_LUT_B97E 16'hB52D
`define CUBE_LUT_B97D 16'hB52B
`define CUBE_LUT_B97C 16'hB528
`define CUBE_LUT_B97B 16'hB525
`define CUBE_LUT_B97A 16'hB522
`define CUBE_LUT_B979 16'hB51F
`define CUBE_LUT_B978 16'hB51C
`define CUBE_LUT_B977 16'hB51A
`define CUBE_LUT_B976 16'hB517
`define CUBE_LUT_B975 16'hB514
`define CUBE_LUT_B974 16'hB511
`define CUBE_LUT_B973 16'hB50E
`define CUBE_LUT_B972 16'hB50C
`define CUBE_LUT_B971 16'hB509
`define CUBE_LUT_B970 16'hB506
`define CUBE_LUT_B96F 16'hB503
`define CUBE_LUT_B96E 16'hB501
`define CUBE_LUT_B96D 16'hB4FE
`define CUBE_LUT_B96C 16'hB4FB
`define CUBE_LUT_B96B 16'hB4F8
`define CUBE_LUT_B96A 16'hB4F6
`define CUBE_LUT_B969 16'hB4F3
`define CUBE_LUT_B968 16'hB4F0
`define CUBE_LUT_B967 16'hB4ED
`define CUBE_LUT_B966 16'hB4EB
`define CUBE_LUT_B965 16'hB4E8
`define CUBE_LUT_B964 16'hB4E5
`define CUBE_LUT_B963 16'hB4E2
`define CUBE_LUT_B962 16'hB4E0
`define CUBE_LUT_B961 16'hB4DD
`define CUBE_LUT_B960 16'hB4DA
`define CUBE_LUT_B95F 16'hB4D8
`define CUBE_LUT_B95E 16'hB4D5
`define CUBE_LUT_B95D 16'hB4D2
`define CUBE_LUT_B95C 16'hB4CF
`define CUBE_LUT_B95B 16'hB4CD
`define CUBE_LUT_B95A 16'hB4CA
`define CUBE_LUT_B959 16'hB4C7
`define CUBE_LUT_B958 16'hB4C5
`define CUBE_LUT_B957 16'hB4C2
`define CUBE_LUT_B956 16'hB4BF
`define CUBE_LUT_B955 16'hB4BD
`define CUBE_LUT_B954 16'hB4BA
`define CUBE_LUT_B953 16'hB4B7
`define CUBE_LUT_B952 16'hB4B5
`define CUBE_LUT_B951 16'hB4B2
`define CUBE_LUT_B950 16'hB4AF
`define CUBE_LUT_B94F 16'hB4AD
`define CUBE_LUT_B94E 16'hB4AA
`define CUBE_LUT_B94D 16'hB4A8
`define CUBE_LUT_B94C 16'hB4A5
`define CUBE_LUT_B94B 16'hB4A2
`define CUBE_LUT_B94A 16'hB4A0
`define CUBE_LUT_B949 16'hB49D
`define CUBE_LUT_B948 16'hB49A
`define CUBE_LUT_B947 16'hB498
`define CUBE_LUT_B946 16'hB495
`define CUBE_LUT_B945 16'hB493
`define CUBE_LUT_B944 16'hB490
`define CUBE_LUT_B943 16'hB48D
`define CUBE_LUT_B942 16'hB48B
`define CUBE_LUT_B941 16'hB488
`define CUBE_LUT_B940 16'hB486
`define CUBE_LUT_B93F 16'hB483
`define CUBE_LUT_B93E 16'hB480
`define CUBE_LUT_B93D 16'hB47E
`define CUBE_LUT_B93C 16'hB47B
`define CUBE_LUT_B93B 16'hB479
`define CUBE_LUT_B93A 16'hB476
`define CUBE_LUT_B939 16'hB474
`define CUBE_LUT_B938 16'hB471
`define CUBE_LUT_B937 16'hB46F
`define CUBE_LUT_B936 16'hB46C
`define CUBE_LUT_B935 16'hB469
`define CUBE_LUT_B934 16'hB467
`define CUBE_LUT_B933 16'hB464
`define CUBE_LUT_B932 16'hB462
`define CUBE_LUT_B931 16'hB45F
`define CUBE_LUT_B930 16'hB45D
`define CUBE_LUT_B92F 16'hB45A
`define CUBE_LUT_B92E 16'hB458
`define CUBE_LUT_B92D 16'hB455
`define CUBE_LUT_B92C 16'hB453
`define CUBE_LUT_B92B 16'hB450
`define CUBE_LUT_B92A 16'hB44E
`define CUBE_LUT_B929 16'hB44B
`define CUBE_LUT_B928 16'hB449
`define CUBE_LUT_B927 16'hB446
`define CUBE_LUT_B926 16'hB444
`define CUBE_LUT_B925 16'hB441
`define CUBE_LUT_B924 16'hB43F
`define CUBE_LUT_B923 16'hB43C
`define CUBE_LUT_B922 16'hB43A
`define CUBE_LUT_B921 16'hB437
`define CUBE_LUT_B920 16'hB435
`define CUBE_LUT_B91F 16'hB432
`define CUBE_LUT_B91E 16'hB430
`define CUBE_LUT_B91D 16'hB42E
`define CUBE_LUT_B91C 16'hB42B
`define CUBE_LUT_B91B 16'hB429
`define CUBE_LUT_B91A 16'hB426
`define CUBE_LUT_B919 16'hB424
`define CUBE_LUT_B918 16'hB421
`define CUBE_LUT_B917 16'hB41F
`define CUBE_LUT_B916 16'hB41C
`define CUBE_LUT_B915 16'hB41A
`define CUBE_LUT_B914 16'hB418
`define CUBE_LUT_B913 16'hB415
`define CUBE_LUT_B912 16'hB413
`define CUBE_LUT_B911 16'hB410
`define CUBE_LUT_B910 16'hB40E
`define CUBE_LUT_B90F 16'hB40C
`define CUBE_LUT_B90E 16'hB409
`define CUBE_LUT_B90D 16'hB407
`define CUBE_LUT_B90C 16'hB404
`define CUBE_LUT_B90B 16'hB402
`define CUBE_LUT_B90A 16'hB3FF
`define CUBE_LUT_B909 16'hB3FA
`define CUBE_LUT_B908 16'hB3F6
`define CUBE_LUT_B907 16'hB3F1
`define CUBE_LUT_B906 16'hB3EC
`define CUBE_LUT_B905 16'hB3E8
`define CUBE_LUT_B904 16'hB3E3
`define CUBE_LUT_B903 16'hB3DE
`define CUBE_LUT_B902 16'hB3D9
`define CUBE_LUT_B901 16'hB3D5
`define CUBE_LUT_B900 16'hB3D0
`define CUBE_LUT_B8FF 16'hB3CB
`define CUBE_LUT_B8FE 16'hB3C7
`define CUBE_LUT_B8FD 16'hB3C2
`define CUBE_LUT_B8FC 16'hB3BD
`define CUBE_LUT_B8FB 16'hB3B9
`define CUBE_LUT_B8FA 16'hB3B4
`define CUBE_LUT_B8F9 16'hB3AF
`define CUBE_LUT_B8F8 16'hB3AB
`define CUBE_LUT_B8F7 16'hB3A6
`define CUBE_LUT_B8F6 16'hB3A1
`define CUBE_LUT_B8F5 16'hB39D
`define CUBE_LUT_B8F4 16'hB398
`define CUBE_LUT_B8F3 16'hB394
`define CUBE_LUT_B8F2 16'hB38F
`define CUBE_LUT_B8F1 16'hB38B
`define CUBE_LUT_B8F0 16'hB386
`define CUBE_LUT_B8EF 16'hB381
`define CUBE_LUT_B8EE 16'hB37D
`define CUBE_LUT_B8ED 16'hB378
`define CUBE_LUT_B8EC 16'hB374
`define CUBE_LUT_B8EB 16'hB36F
`define CUBE_LUT_B8EA 16'hB36B
`define CUBE_LUT_B8E9 16'hB366
`define CUBE_LUT_B8E8 16'hB362
`define CUBE_LUT_B8E7 16'hB35D
`define CUBE_LUT_B8E6 16'hB359
`define CUBE_LUT_B8E5 16'hB354
`define CUBE_LUT_B8E4 16'hB350
`define CUBE_LUT_B8E3 16'hB34B
`define CUBE_LUT_B8E2 16'hB347
`define CUBE_LUT_B8E1 16'hB342
`define CUBE_LUT_B8E0 16'hB33E
`define CUBE_LUT_B8DF 16'hB339
`define CUBE_LUT_B8DE 16'hB335
`define CUBE_LUT_B8DD 16'hB330
`define CUBE_LUT_B8DC 16'hB32C
`define CUBE_LUT_B8DB 16'hB328
`define CUBE_LUT_B8DA 16'hB323
`define CUBE_LUT_B8D9 16'hB31F
`define CUBE_LUT_B8D8 16'hB31A
`define CUBE_LUT_B8D7 16'hB316
`define CUBE_LUT_B8D6 16'hB312
`define CUBE_LUT_B8D5 16'hB30D
`define CUBE_LUT_B8D4 16'hB309
`define CUBE_LUT_B8D3 16'hB304
`define CUBE_LUT_B8D2 16'hB300
`define CUBE_LUT_B8D1 16'hB2FC
`define CUBE_LUT_B8D0 16'hB2F7
`define CUBE_LUT_B8CF 16'hB2F3
`define CUBE_LUT_B8CE 16'hB2EF
`define CUBE_LUT_B8CD 16'hB2EA
`define CUBE_LUT_B8CC 16'hB2E6
`define CUBE_LUT_B8CB 16'hB2E2
`define CUBE_LUT_B8CA 16'hB2DD
`define CUBE_LUT_B8C9 16'hB2D9
`define CUBE_LUT_B8C8 16'hB2D5
`define CUBE_LUT_B8C7 16'hB2D1
`define CUBE_LUT_B8C6 16'hB2CC
`define CUBE_LUT_B8C5 16'hB2C8
`define CUBE_LUT_B8C4 16'hB2C4
`define CUBE_LUT_B8C3 16'hB2BF
`define CUBE_LUT_B8C2 16'hB2BB
`define CUBE_LUT_B8C1 16'hB2B7
`define CUBE_LUT_B8C0 16'hB2B3
`define CUBE_LUT_B8BF 16'hB2AF
`define CUBE_LUT_B8BE 16'hB2AA
`define CUBE_LUT_B8BD 16'hB2A6
`define CUBE_LUT_B8BC 16'hB2A2
`define CUBE_LUT_B8BB 16'hB29E
`define CUBE_LUT_B8BA 16'hB299
`define CUBE_LUT_B8B9 16'hB295
`define CUBE_LUT_B8B8 16'hB291
`define CUBE_LUT_B8B7 16'hB28D
`define CUBE_LUT_B8B6 16'hB289
`define CUBE_LUT_B8B5 16'hB285
`define CUBE_LUT_B8B4 16'hB280
`define CUBE_LUT_B8B3 16'hB27C
`define CUBE_LUT_B8B2 16'hB278
`define CUBE_LUT_B8B1 16'hB274
`define CUBE_LUT_B8B0 16'hB270
`define CUBE_LUT_B8AF 16'hB26C
`define CUBE_LUT_B8AE 16'hB268
`define CUBE_LUT_B8AD 16'hB264
`define CUBE_LUT_B8AC 16'hB260
`define CUBE_LUT_B8AB 16'hB25B
`define CUBE_LUT_B8AA 16'hB257
`define CUBE_LUT_B8A9 16'hB253
`define CUBE_LUT_B8A8 16'hB24F
`define CUBE_LUT_B8A7 16'hB24B
`define CUBE_LUT_B8A6 16'hB247
`define CUBE_LUT_B8A5 16'hB243
`define CUBE_LUT_B8A4 16'hB23F
`define CUBE_LUT_B8A3 16'hB23B
`define CUBE_LUT_B8A2 16'hB237
`define CUBE_LUT_B8A1 16'hB233
`define CUBE_LUT_B8A0 16'hB22F
`define CUBE_LUT_B89F 16'hB22B
`define CUBE_LUT_B89E 16'hB227
`define CUBE_LUT_B89D 16'hB223
`define CUBE_LUT_B89C 16'hB21F
`define CUBE_LUT_B89B 16'hB21B
`define CUBE_LUT_B89A 16'hB217
`define CUBE_LUT_B899 16'hB213
`define CUBE_LUT_B898 16'hB20F
`define CUBE_LUT_B897 16'hB20B
`define CUBE_LUT_B896 16'hB207
`define CUBE_LUT_B895 16'hB203
`define CUBE_LUT_B894 16'hB1FF
`define CUBE_LUT_B893 16'hB1FB
`define CUBE_LUT_B892 16'hB1F7
`define CUBE_LUT_B891 16'hB1F4
`define CUBE_LUT_B890 16'hB1F0
`define CUBE_LUT_B88F 16'hB1EC
`define CUBE_LUT_B88E 16'hB1E8
`define CUBE_LUT_B88D 16'hB1E4
`define CUBE_LUT_B88C 16'hB1E0
`define CUBE_LUT_B88B 16'hB1DC
`define CUBE_LUT_B88A 16'hB1D8
`define CUBE_LUT_B889 16'hB1D4
`define CUBE_LUT_B888 16'hB1D1
`define CUBE_LUT_B887 16'hB1CD
`define CUBE_LUT_B886 16'hB1C9
`define CUBE_LUT_B885 16'hB1C5
`define CUBE_LUT_B884 16'hB1C1
`define CUBE_LUT_B883 16'hB1BD
`define CUBE_LUT_B882 16'hB1BA
`define CUBE_LUT_B881 16'hB1B6
`define CUBE_LUT_B880 16'hB1B2
`define CUBE_LUT_B87F 16'hB1AE
`define CUBE_LUT_B87E 16'hB1AA
`define CUBE_LUT_B87D 16'hB1A7
`define CUBE_LUT_B87C 16'hB1A3
`define CUBE_LUT_B87B 16'hB19F
`define CUBE_LUT_B87A 16'hB19B
`define CUBE_LUT_B879 16'hB198
`define CUBE_LUT_B878 16'hB194
`define CUBE_LUT_B877 16'hB190
`define CUBE_LUT_B876 16'hB18C
`define CUBE_LUT_B875 16'hB189
`define CUBE_LUT_B874 16'hB185
`define CUBE_LUT_B873 16'hB181
`define CUBE_LUT_B872 16'hB17D
`define CUBE_LUT_B871 16'hB17A
`define CUBE_LUT_B870 16'hB176
`define CUBE_LUT_B86F 16'hB172
`define CUBE_LUT_B86E 16'hB16F
`define CUBE_LUT_B86D 16'hB16B
`define CUBE_LUT_B86C 16'hB167
`define CUBE_LUT_B86B 16'hB164
`define CUBE_LUT_B86A 16'hB160
`define CUBE_LUT_B869 16'hB15C
`define CUBE_LUT_B868 16'hB159
`define CUBE_LUT_B867 16'hB155
`define CUBE_LUT_B866 16'hB151
`define CUBE_LUT_B865 16'hB14E
`define CUBE_LUT_B864 16'hB14A
`define CUBE_LUT_B863 16'hB147
`define CUBE_LUT_B862 16'hB143
`define CUBE_LUT_B861 16'hB13F
`define CUBE_LUT_B860 16'hB13C
`define CUBE_LUT_B85F 16'hB138
`define CUBE_LUT_B85E 16'hB135
`define CUBE_LUT_B85D 16'hB131
`define CUBE_LUT_B85C 16'hB12E
`define CUBE_LUT_B85B 16'hB12A
`define CUBE_LUT_B85A 16'hB126
`define CUBE_LUT_B859 16'hB123
`define CUBE_LUT_B858 16'hB11F
`define CUBE_LUT_B857 16'hB11C
`define CUBE_LUT_B856 16'hB118
`define CUBE_LUT_B855 16'hB115
`define CUBE_LUT_B854 16'hB111
`define CUBE_LUT_B853 16'hB10E
`define CUBE_LUT_B852 16'hB10A
`define CUBE_LUT_B851 16'hB107
`define CUBE_LUT_B850 16'hB103
`define CUBE_LUT_B84F 16'hB100
`define CUBE_LUT_B84E 16'hB0FC
`define CUBE_LUT_B84D 16'hB0F9
`define CUBE_LUT_B84C 16'hB0F5
`define CUBE_LUT_B84B 16'hB0F2
`define CUBE_LUT_B84A 16'hB0EE
`define CUBE_LUT_B849 16'hB0EB
`define CUBE_LUT_B848 16'hB0E8
`define CUBE_LUT_B847 16'hB0E4
`define CUBE_LUT_B846 16'hB0E1
`define CUBE_LUT_B845 16'hB0DD
`define CUBE_LUT_B844 16'hB0DA
`define CUBE_LUT_B843 16'hB0D6
`define CUBE_LUT_B842 16'hB0D3
`define CUBE_LUT_B841 16'hB0D0
`define CUBE_LUT_B840 16'hB0CC
`define CUBE_LUT_B83F 16'hB0C9
`define CUBE_LUT_B83E 16'hB0C5
`define CUBE_LUT_B83D 16'hB0C2
`define CUBE_LUT_B83C 16'hB0BF
`define CUBE_LUT_B83B 16'hB0BB
`define CUBE_LUT_B83A 16'hB0B8
`define CUBE_LUT_B839 16'hB0B5
`define CUBE_LUT_B838 16'hB0B1
`define CUBE_LUT_B837 16'hB0AE
`define CUBE_LUT_B836 16'hB0AB
`define CUBE_LUT_B835 16'hB0A7
`define CUBE_LUT_B834 16'hB0A4
`define CUBE_LUT_B833 16'hB0A1
`define CUBE_LUT_B832 16'hB09D
`define CUBE_LUT_B831 16'hB09A
`define CUBE_LUT_B830 16'hB097
`define CUBE_LUT_B82F 16'hB094
`define CUBE_LUT_B82E 16'hB090
`define CUBE_LUT_B82D 16'hB08D
`define CUBE_LUT_B82C 16'hB08A
`define CUBE_LUT_B82B 16'hB086
`define CUBE_LUT_B82A 16'hB083
`define CUBE_LUT_B829 16'hB080
`define CUBE_LUT_B828 16'hB07D
`define CUBE_LUT_B827 16'hB07A
`define CUBE_LUT_B826 16'hB076
`define CUBE_LUT_B825 16'hB073
`define CUBE_LUT_B824 16'hB070
`define CUBE_LUT_B823 16'hB06D
`define CUBE_LUT_B822 16'hB069
`define CUBE_LUT_B821 16'hB066
`define CUBE_LUT_B820 16'hB063
`define CUBE_LUT_B81F 16'hB060
`define CUBE_LUT_B81E 16'hB05D
`define CUBE_LUT_B81D 16'hB059
`define CUBE_LUT_B81C 16'hB056
`define CUBE_LUT_B81B 16'hB053
`define CUBE_LUT_B81A 16'hB050
`define CUBE_LUT_B819 16'hB04D
`define CUBE_LUT_B818 16'hB04A
`define CUBE_LUT_B817 16'hB047
`define CUBE_LUT_B816 16'hB043
`define CUBE_LUT_B815 16'hB040
`define CUBE_LUT_B814 16'hB03D
`define CUBE_LUT_B813 16'hB03A
`define CUBE_LUT_B812 16'hB037
`define CUBE_LUT_B811 16'hB034
`define CUBE_LUT_B810 16'hB031
`define CUBE_LUT_B80F 16'hB02E
`define CUBE_LUT_B80E 16'hB02B
`define CUBE_LUT_B80D 16'hB027
`define CUBE_LUT_B80C 16'hB024
`define CUBE_LUT_B80B 16'hB021
`define CUBE_LUT_B80A 16'hB01E
`define CUBE_LUT_B809 16'hB01B
`define CUBE_LUT_B808 16'hB018
`define CUBE_LUT_B807 16'hB015
`define CUBE_LUT_B806 16'hB012
`define CUBE_LUT_B805 16'hB00F
`define CUBE_LUT_B804 16'hB00C
`define CUBE_LUT_B803 16'hB009
`define CUBE_LUT_B802 16'hB006
`define CUBE_LUT_B801 16'hB003
`define CUBE_LUT_B800 16'hB000
`define CUBE_LUT_B7FF 16'hAFFD
`define CUBE_LUT_B7FE 16'hAFFA
`define CUBE_LUT_B7FD 16'hAFF7
`define CUBE_LUT_B7FC 16'hAFF4
`define CUBE_LUT_B7FB 16'hAFF1
`define CUBE_LUT_B7FA 16'hAFEE
`define CUBE_LUT_B7F9 16'hAFEB
`define CUBE_LUT_B7F8 16'hAFE8
`define CUBE_LUT_B7F7 16'hAFE5
`define CUBE_LUT_B7F6 16'hAFE2
`define CUBE_LUT_B7F5 16'hAFDF
`define CUBE_LUT_B7F4 16'hAFDC
`define CUBE_LUT_B7F3 16'hAFD9
`define CUBE_LUT_B7F2 16'hAFD6
`define CUBE_LUT_B7F1 16'hAFD3
`define CUBE_LUT_B7F0 16'hAFD0
`define CUBE_LUT_B7EF 16'hAFCD
`define CUBE_LUT_B7EE 16'hAFCA
`define CUBE_LUT_B7ED 16'hAFC8
`define CUBE_LUT_B7EC 16'hAFC5
`define CUBE_LUT_B7EB 16'hAFC2
`define CUBE_LUT_B7EA 16'hAFBF
`define CUBE_LUT_B7E9 16'hAFBC
`define CUBE_LUT_B7E8 16'hAFB9
`define CUBE_LUT_B7E7 16'hAFB6
`define CUBE_LUT_B7E6 16'hAFB3
`define CUBE_LUT_B7E5 16'hAFB0
`define CUBE_LUT_B7E4 16'hAFAD
`define CUBE_LUT_B7E3 16'hAFAA
`define CUBE_LUT_B7E2 16'hAFA7
`define CUBE_LUT_B7E1 16'hAFA4
`define CUBE_LUT_B7E0 16'hAFA1
`define CUBE_LUT_B7DF 16'hAF9F
`define CUBE_LUT_B7DE 16'hAF9C
`define CUBE_LUT_B7DD 16'hAF99
`define CUBE_LUT_B7DC 16'hAF96
`define CUBE_LUT_B7DB 16'hAF93
`define CUBE_LUT_B7DA 16'hAF90
`define CUBE_LUT_B7D9 16'hAF8D
`define CUBE_LUT_B7D8 16'hAF8A
`define CUBE_LUT_B7D7 16'hAF87
`define CUBE_LUT_B7D6 16'hAF85
`define CUBE_LUT_B7D5 16'hAF82
`define CUBE_LUT_B7D4 16'hAF7F
`define CUBE_LUT_B7D3 16'hAF7C
`define CUBE_LUT_B7D2 16'hAF79
`define CUBE_LUT_B7D1 16'hAF76
`define CUBE_LUT_B7D0 16'hAF73
`define CUBE_LUT_B7CF 16'hAF70
`define CUBE_LUT_B7CE 16'hAF6E
`define CUBE_LUT_B7CD 16'hAF6B
`define CUBE_LUT_B7CC 16'hAF68
`define CUBE_LUT_B7CB 16'hAF65
`define CUBE_LUT_B7CA 16'hAF62
`define CUBE_LUT_B7C9 16'hAF5F
`define CUBE_LUT_B7C8 16'hAF5D
`define CUBE_LUT_B7C7 16'hAF5A
`define CUBE_LUT_B7C6 16'hAF57
`define CUBE_LUT_B7C5 16'hAF54
`define CUBE_LUT_B7C4 16'hAF51
`define CUBE_LUT_B7C3 16'hAF4E
`define CUBE_LUT_B7C2 16'hAF4C
`define CUBE_LUT_B7C1 16'hAF49
`define CUBE_LUT_B7C0 16'hAF46
`define CUBE_LUT_B7BF 16'hAF43
`define CUBE_LUT_B7BE 16'hAF40
`define CUBE_LUT_B7BD 16'hAF3E
`define CUBE_LUT_B7BC 16'hAF3B
`define CUBE_LUT_B7BB 16'hAF38
`define CUBE_LUT_B7BA 16'hAF35
`define CUBE_LUT_B7B9 16'hAF32
`define CUBE_LUT_B7B8 16'hAF30
`define CUBE_LUT_B7B7 16'hAF2D
`define CUBE_LUT_B7B6 16'hAF2A
`define CUBE_LUT_B7B5 16'hAF27
`define CUBE_LUT_B7B4 16'hAF24
`define CUBE_LUT_B7B3 16'hAF22
`define CUBE_LUT_B7B2 16'hAF1F
`define CUBE_LUT_B7B1 16'hAF1C
`define CUBE_LUT_B7B0 16'hAF19
`define CUBE_LUT_B7AF 16'hAF16
`define CUBE_LUT_B7AE 16'hAF14
`define CUBE_LUT_B7AD 16'hAF11
`define CUBE_LUT_B7AC 16'hAF0E
`define CUBE_LUT_B7AB 16'hAF0B
`define CUBE_LUT_B7AA 16'hAF09
`define CUBE_LUT_B7A9 16'hAF06
`define CUBE_LUT_B7A8 16'hAF03
`define CUBE_LUT_B7A7 16'hAF00
`define CUBE_LUT_B7A6 16'hAEFE
`define CUBE_LUT_B7A5 16'hAEFB
`define CUBE_LUT_B7A4 16'hAEF8
`define CUBE_LUT_B7A3 16'hAEF5
`define CUBE_LUT_B7A2 16'hAEF3
`define CUBE_LUT_B7A1 16'hAEF0
`define CUBE_LUT_B7A0 16'hAEED
`define CUBE_LUT_B79F 16'hAEEB
`define CUBE_LUT_B79E 16'hAEE8
`define CUBE_LUT_B79D 16'hAEE5
`define CUBE_LUT_B79C 16'hAEE2
`define CUBE_LUT_B79B 16'hAEE0
`define CUBE_LUT_B79A 16'hAEDD
`define CUBE_LUT_B799 16'hAEDA
`define CUBE_LUT_B798 16'hAED8
`define CUBE_LUT_B797 16'hAED5
`define CUBE_LUT_B796 16'hAED2
`define CUBE_LUT_B795 16'hAECF
`define CUBE_LUT_B794 16'hAECD
`define CUBE_LUT_B793 16'hAECA
`define CUBE_LUT_B792 16'hAEC7
`define CUBE_LUT_B791 16'hAEC5
`define CUBE_LUT_B790 16'hAEC2
`define CUBE_LUT_B78F 16'hAEBF
`define CUBE_LUT_B78E 16'hAEBD
`define CUBE_LUT_B78D 16'hAEBA
`define CUBE_LUT_B78C 16'hAEB7
`define CUBE_LUT_B78B 16'hAEB5
`define CUBE_LUT_B78A 16'hAEB2
`define CUBE_LUT_B789 16'hAEAF
`define CUBE_LUT_B788 16'hAEAD
`define CUBE_LUT_B787 16'hAEAA
`define CUBE_LUT_B786 16'hAEA7
`define CUBE_LUT_B785 16'hAEA5
`define CUBE_LUT_B784 16'hAEA2
`define CUBE_LUT_B783 16'hAE9F
`define CUBE_LUT_B782 16'hAE9D
`define CUBE_LUT_B781 16'hAE9A
`define CUBE_LUT_B780 16'hAE98
`define CUBE_LUT_B77F 16'hAE95
`define CUBE_LUT_B77E 16'hAE92
`define CUBE_LUT_B77D 16'hAE90
`define CUBE_LUT_B77C 16'hAE8D
`define CUBE_LUT_B77B 16'hAE8A
`define CUBE_LUT_B77A 16'hAE88
`define CUBE_LUT_B779 16'hAE85
`define CUBE_LUT_B778 16'hAE82
`define CUBE_LUT_B777 16'hAE80
`define CUBE_LUT_B776 16'hAE7D
`define CUBE_LUT_B775 16'hAE7B
`define CUBE_LUT_B774 16'hAE78
`define CUBE_LUT_B773 16'hAE75
`define CUBE_LUT_B772 16'hAE73
`define CUBE_LUT_B771 16'hAE70
`define CUBE_LUT_B770 16'hAE6E
`define CUBE_LUT_B76F 16'hAE6B
`define CUBE_LUT_B76E 16'hAE68
`define CUBE_LUT_B76D 16'hAE66
`define CUBE_LUT_B76C 16'hAE63
`define CUBE_LUT_B76B 16'hAE61
`define CUBE_LUT_B76A 16'hAE5E
`define CUBE_LUT_B769 16'hAE5C
`define CUBE_LUT_B768 16'hAE59
`define CUBE_LUT_B767 16'hAE56
`define CUBE_LUT_B766 16'hAE54
`define CUBE_LUT_B765 16'hAE51
`define CUBE_LUT_B764 16'hAE4F
`define CUBE_LUT_B763 16'hAE4C
`define CUBE_LUT_B762 16'hAE4A
`define CUBE_LUT_B761 16'hAE47
`define CUBE_LUT_B760 16'hAE45
`define CUBE_LUT_B75F 16'hAE42
`define CUBE_LUT_B75E 16'hAE3F
`define CUBE_LUT_B75D 16'hAE3D
`define CUBE_LUT_B75C 16'hAE3A
`define CUBE_LUT_B75B 16'hAE38
`define CUBE_LUT_B75A 16'hAE35
`define CUBE_LUT_B759 16'hAE33
`define CUBE_LUT_B758 16'hAE30
`define CUBE_LUT_B757 16'hAE2E
`define CUBE_LUT_B756 16'hAE2B
`define CUBE_LUT_B755 16'hAE29
`define CUBE_LUT_B754 16'hAE26
`define CUBE_LUT_B753 16'hAE24
`define CUBE_LUT_B752 16'hAE21
`define CUBE_LUT_B751 16'hAE1F
`define CUBE_LUT_B750 16'hAE1C
`define CUBE_LUT_B74F 16'hAE1A
`define CUBE_LUT_B74E 16'hAE17
`define CUBE_LUT_B74D 16'hAE15
`define CUBE_LUT_B74C 16'hAE12
`define CUBE_LUT_B74B 16'hAE10
`define CUBE_LUT_B74A 16'hAE0D
`define CUBE_LUT_B749 16'hAE0B
`define CUBE_LUT_B748 16'hAE08
`define CUBE_LUT_B747 16'hAE06
`define CUBE_LUT_B746 16'hAE03
`define CUBE_LUT_B745 16'hAE01
`define CUBE_LUT_B744 16'hADFE
`define CUBE_LUT_B743 16'hADFC
`define CUBE_LUT_B742 16'hADF9
`define CUBE_LUT_B741 16'hADF7
`define CUBE_LUT_B740 16'hADF4
`define CUBE_LUT_B73F 16'hADF2
`define CUBE_LUT_B73E 16'hADEF
`define CUBE_LUT_B73D 16'hADED
`define CUBE_LUT_B73C 16'hADEA
`define CUBE_LUT_B73B 16'hADE8
`define CUBE_LUT_B73A 16'hADE6
`define CUBE_LUT_B739 16'hADE3
`define CUBE_LUT_B738 16'hADE1
`define CUBE_LUT_B737 16'hADDE
`define CUBE_LUT_B736 16'hADDC
`define CUBE_LUT_B735 16'hADD9
`define CUBE_LUT_B734 16'hADD7
`define CUBE_LUT_B733 16'hADD5
`define CUBE_LUT_B732 16'hADD2
`define CUBE_LUT_B731 16'hADD0
`define CUBE_LUT_B730 16'hADCD
`define CUBE_LUT_B72F 16'hADCB
`define CUBE_LUT_B72E 16'hADC8
`define CUBE_LUT_B72D 16'hADC6
`define CUBE_LUT_B72C 16'hADC4
`define CUBE_LUT_B72B 16'hADC1
`define CUBE_LUT_B72A 16'hADBF
`define CUBE_LUT_B729 16'hADBC
`define CUBE_LUT_B728 16'hADBA
`define CUBE_LUT_B727 16'hADB8
`define CUBE_LUT_B726 16'hADB5
`define CUBE_LUT_B725 16'hADB3
`define CUBE_LUT_B724 16'hADB0
`define CUBE_LUT_B723 16'hADAE
`define CUBE_LUT_B722 16'hADAC
`define CUBE_LUT_B721 16'hADA9
`define CUBE_LUT_B720 16'hADA7
`define CUBE_LUT_B71F 16'hADA4
`define CUBE_LUT_B71E 16'hADA2
`define CUBE_LUT_B71D 16'hADA0
`define CUBE_LUT_B71C 16'hAD9D
`define CUBE_LUT_B71B 16'hAD9B
`define CUBE_LUT_B71A 16'hAD99
`define CUBE_LUT_B719 16'hAD96
`define CUBE_LUT_B718 16'hAD94
`define CUBE_LUT_B717 16'hAD92
`define CUBE_LUT_B716 16'hAD8F
`define CUBE_LUT_B715 16'hAD8D
`define CUBE_LUT_B714 16'hAD8A
`define CUBE_LUT_B713 16'hAD88
`define CUBE_LUT_B712 16'hAD86
`define CUBE_LUT_B711 16'hAD83
`define CUBE_LUT_B710 16'hAD81
`define CUBE_LUT_B70F 16'hAD7F
`define CUBE_LUT_B70E 16'hAD7C
`define CUBE_LUT_B70D 16'hAD7A
`define CUBE_LUT_B70C 16'hAD78
`define CUBE_LUT_B70B 16'hAD75
`define CUBE_LUT_B70A 16'hAD73
`define CUBE_LUT_B709 16'hAD71
`define CUBE_LUT_B708 16'hAD6E
`define CUBE_LUT_B707 16'hAD6C
`define CUBE_LUT_B706 16'hAD6A
`define CUBE_LUT_B705 16'hAD68
`define CUBE_LUT_B704 16'hAD65
`define CUBE_LUT_B703 16'hAD63
`define CUBE_LUT_B702 16'hAD61
`define CUBE_LUT_B701 16'hAD5E
`define CUBE_LUT_B700 16'hAD5C
`define CUBE_LUT_B6FF 16'hAD5A
`define CUBE_LUT_B6FE 16'hAD57
`define CUBE_LUT_B6FD 16'hAD55
`define CUBE_LUT_B6FC 16'hAD53
`define CUBE_LUT_B6FB 16'hAD51
`define CUBE_LUT_B6FA 16'hAD4E
`define CUBE_LUT_B6F9 16'hAD4C
`define CUBE_LUT_B6F8 16'hAD4A
`define CUBE_LUT_B6F7 16'hAD47
`define CUBE_LUT_B6F6 16'hAD45
`define CUBE_LUT_B6F5 16'hAD43
`define CUBE_LUT_B6F4 16'hAD41
`define CUBE_LUT_B6F3 16'hAD3E
`define CUBE_LUT_B6F2 16'hAD3C
`define CUBE_LUT_B6F1 16'hAD3A
`define CUBE_LUT_B6F0 16'hAD38
`define CUBE_LUT_B6EF 16'hAD35
`define CUBE_LUT_B6EE 16'hAD33
`define CUBE_LUT_B6ED 16'hAD31
`define CUBE_LUT_B6EC 16'hAD2F
`define CUBE_LUT_B6EB 16'hAD2C
`define CUBE_LUT_B6EA 16'hAD2A
`define CUBE_LUT_B6E9 16'hAD28
`define CUBE_LUT_B6E8 16'hAD26
`define CUBE_LUT_B6E7 16'hAD23
`define CUBE_LUT_B6E6 16'hAD21
`define CUBE_LUT_B6E5 16'hAD1F
`define CUBE_LUT_B6E4 16'hAD1D
`define CUBE_LUT_B6E3 16'hAD1A
`define CUBE_LUT_B6E2 16'hAD18
`define CUBE_LUT_B6E1 16'hAD16
`define CUBE_LUT_B6E0 16'hAD14
`define CUBE_LUT_B6DF 16'hAD12
`define CUBE_LUT_B6DE 16'hAD0F
`define CUBE_LUT_B6DD 16'hAD0D
`define CUBE_LUT_B6DC 16'hAD0B
`define CUBE_LUT_B6DB 16'hAD09
`define CUBE_LUT_B6DA 16'hAD07
`define CUBE_LUT_B6D9 16'hAD04
`define CUBE_LUT_B6D8 16'hAD02
`define CUBE_LUT_B6D7 16'hAD00
`define CUBE_LUT_B6D6 16'hACFE
`define CUBE_LUT_B6D5 16'hACFC
`define CUBE_LUT_B6D4 16'hACF9
`define CUBE_LUT_B6D3 16'hACF7
`define CUBE_LUT_B6D2 16'hACF5
`define CUBE_LUT_B6D1 16'hACF3
`define CUBE_LUT_B6D0 16'hACF1
`define CUBE_LUT_B6CF 16'hACEF
`define CUBE_LUT_B6CE 16'hACEC
`define CUBE_LUT_B6CD 16'hACEA
`define CUBE_LUT_B6CC 16'hACE8
`define CUBE_LUT_B6CB 16'hACE6
`define CUBE_LUT_B6CA 16'hACE4
`define CUBE_LUT_B6C9 16'hACE2
`define CUBE_LUT_B6C8 16'hACDF
`define CUBE_LUT_B6C7 16'hACDD
`define CUBE_LUT_B6C6 16'hACDB
`define CUBE_LUT_B6C5 16'hACD9
`define CUBE_LUT_B6C4 16'hACD7
`define CUBE_LUT_B6C3 16'hACD5
`define CUBE_LUT_B6C2 16'hACD2
`define CUBE_LUT_B6C1 16'hACD0
`define CUBE_LUT_B6C0 16'hACCE
`define CUBE_LUT_B6BF 16'hACCC
`define CUBE_LUT_B6BE 16'hACCA
`define CUBE_LUT_B6BD 16'hACC8
`define CUBE_LUT_B6BC 16'hACC6
`define CUBE_LUT_B6BB 16'hACC4
`define CUBE_LUT_B6BA 16'hACC1
`define CUBE_LUT_B6B9 16'hACBF
`define CUBE_LUT_B6B8 16'hACBD
`define CUBE_LUT_B6B7 16'hACBB
`define CUBE_LUT_B6B6 16'hACB9
`define CUBE_LUT_B6B5 16'hACB7
`define CUBE_LUT_B6B4 16'hACB5
`define CUBE_LUT_B6B3 16'hACB3
`define CUBE_LUT_B6B2 16'hACB1
`define CUBE_LUT_B6B1 16'hACAE
`define CUBE_LUT_B6B0 16'hACAC
`define CUBE_LUT_B6AF 16'hACAA
`define CUBE_LUT_B6AE 16'hACA8
`define CUBE_LUT_B6AD 16'hACA6
`define CUBE_LUT_B6AC 16'hACA4
`define CUBE_LUT_B6AB 16'hACA2
`define CUBE_LUT_B6AA 16'hACA0
`define CUBE_LUT_B6A9 16'hAC9E
`define CUBE_LUT_B6A8 16'hAC9C
`define CUBE_LUT_B6A7 16'hAC9A
`define CUBE_LUT_B6A6 16'hAC97
`define CUBE_LUT_B6A5 16'hAC95
`define CUBE_LUT_B6A4 16'hAC93
`define CUBE_LUT_B6A3 16'hAC91
`define CUBE_LUT_B6A2 16'hAC8F
`define CUBE_LUT_B6A1 16'hAC8D
`define CUBE_LUT_B6A0 16'hAC8B
`define CUBE_LUT_B69F 16'hAC89
`define CUBE_LUT_B69E 16'hAC87
`define CUBE_LUT_B69D 16'hAC85
`define CUBE_LUT_B69C 16'hAC83
`define CUBE_LUT_B69B 16'hAC81
`define CUBE_LUT_B69A 16'hAC7F
`define CUBE_LUT_B699 16'hAC7D
`define CUBE_LUT_B698 16'hAC7B
`define CUBE_LUT_B697 16'hAC79
`define CUBE_LUT_B696 16'hAC77
`define CUBE_LUT_B695 16'hAC75
`define CUBE_LUT_B694 16'hAC73
`define CUBE_LUT_B693 16'hAC71
`define CUBE_LUT_B692 16'hAC6F
`define CUBE_LUT_B691 16'hAC6D
`define CUBE_LUT_B690 16'hAC6A
`define CUBE_LUT_B68F 16'hAC68
`define CUBE_LUT_B68E 16'hAC66
`define CUBE_LUT_B68D 16'hAC64
`define CUBE_LUT_B68C 16'hAC62
`define CUBE_LUT_B68B 16'hAC60
`define CUBE_LUT_B68A 16'hAC5E
`define CUBE_LUT_B689 16'hAC5C
`define CUBE_LUT_B688 16'hAC5A
`define CUBE_LUT_B687 16'hAC58
`define CUBE_LUT_B686 16'hAC56
`define CUBE_LUT_B685 16'hAC54
`define CUBE_LUT_B684 16'hAC52
`define CUBE_LUT_B683 16'hAC50
`define CUBE_LUT_B682 16'hAC4E
`define CUBE_LUT_B681 16'hAC4C
`define CUBE_LUT_B680 16'hAC4A
`define CUBE_LUT_B67F 16'hAC49
`define CUBE_LUT_B67E 16'hAC47
`define CUBE_LUT_B67D 16'hAC45
`define CUBE_LUT_B67C 16'hAC43
`define CUBE_LUT_B67B 16'hAC41
`define CUBE_LUT_B67A 16'hAC3F
`define CUBE_LUT_B679 16'hAC3D
`define CUBE_LUT_B678 16'hAC3B
`define CUBE_LUT_B677 16'hAC39
`define CUBE_LUT_B676 16'hAC37
`define CUBE_LUT_B675 16'hAC35
`define CUBE_LUT_B674 16'hAC33
`define CUBE_LUT_B673 16'hAC31
`define CUBE_LUT_B672 16'hAC2F
`define CUBE_LUT_B671 16'hAC2D
`define CUBE_LUT_B670 16'hAC2B
`define CUBE_LUT_B66F 16'hAC29
`define CUBE_LUT_B66E 16'hAC27
`define CUBE_LUT_B66D 16'hAC25
`define CUBE_LUT_B66C 16'hAC23
`define CUBE_LUT_B66B 16'hAC21
`define CUBE_LUT_B66A 16'hAC20
`define CUBE_LUT_B669 16'hAC1E
`define CUBE_LUT_B668 16'hAC1C
`define CUBE_LUT_B667 16'hAC1A
`define CUBE_LUT_B666 16'hAC18
`define CUBE_LUT_B665 16'hAC16
`define CUBE_LUT_B664 16'hAC14
`define CUBE_LUT_B663 16'hAC12
`define CUBE_LUT_B662 16'hAC10
`define CUBE_LUT_B661 16'hAC0E
`define CUBE_LUT_B660 16'hAC0C
`define CUBE_LUT_B65F 16'hAC0A
`define CUBE_LUT_B65E 16'hAC09
`define CUBE_LUT_B65D 16'hAC07
`define CUBE_LUT_B65C 16'hAC05
`define CUBE_LUT_B65B 16'hAC03
`define CUBE_LUT_B65A 16'hAC01
`define CUBE_LUT_B659 16'hABFE
`define CUBE_LUT_B658 16'hABFA
`define CUBE_LUT_B657 16'hABF7
`define CUBE_LUT_B656 16'hABF3
`define CUBE_LUT_B655 16'hABEF
`define CUBE_LUT_B654 16'hABEB
`define CUBE_LUT_B653 16'hABE8
`define CUBE_LUT_B652 16'hABE4
`define CUBE_LUT_B651 16'hABE0
`define CUBE_LUT_B650 16'hABDC
`define CUBE_LUT_B64F 16'hABD9
`define CUBE_LUT_B64E 16'hABD5
`define CUBE_LUT_B64D 16'hABD1
`define CUBE_LUT_B64C 16'hABCD
`define CUBE_LUT_B64B 16'hABCA
`define CUBE_LUT_B64A 16'hABC6
`define CUBE_LUT_B649 16'hABC2
`define CUBE_LUT_B648 16'hABBF
`define CUBE_LUT_B647 16'hABBB
`define CUBE_LUT_B646 16'hABB7
`define CUBE_LUT_B645 16'hABB3
`define CUBE_LUT_B644 16'hABB0
`define CUBE_LUT_B643 16'hABAC
`define CUBE_LUT_B642 16'hABA8
`define CUBE_LUT_B641 16'hABA5
`define CUBE_LUT_B640 16'hABA1
`define CUBE_LUT_B63F 16'hAB9D
`define CUBE_LUT_B63E 16'hAB9A
`define CUBE_LUT_B63D 16'hAB96
`define CUBE_LUT_B63C 16'hAB93
`define CUBE_LUT_B63B 16'hAB8F
`define CUBE_LUT_B63A 16'hAB8B
`define CUBE_LUT_B639 16'hAB88
`define CUBE_LUT_B638 16'hAB84
`define CUBE_LUT_B637 16'hAB80
`define CUBE_LUT_B636 16'hAB7D
`define CUBE_LUT_B635 16'hAB79
`define CUBE_LUT_B634 16'hAB76
`define CUBE_LUT_B633 16'hAB72
`define CUBE_LUT_B632 16'hAB6E
`define CUBE_LUT_B631 16'hAB6B
`define CUBE_LUT_B630 16'hAB67
`define CUBE_LUT_B62F 16'hAB64
`define CUBE_LUT_B62E 16'hAB60
`define CUBE_LUT_B62D 16'hAB5C
`define CUBE_LUT_B62C 16'hAB59
`define CUBE_LUT_B62B 16'hAB55
`define CUBE_LUT_B62A 16'hAB52
`define CUBE_LUT_B629 16'hAB4E
`define CUBE_LUT_B628 16'hAB4B
`define CUBE_LUT_B627 16'hAB47
`define CUBE_LUT_B626 16'hAB43
`define CUBE_LUT_B625 16'hAB40
`define CUBE_LUT_B624 16'hAB3C
`define CUBE_LUT_B623 16'hAB39
`define CUBE_LUT_B622 16'hAB35
`define CUBE_LUT_B621 16'hAB32
`define CUBE_LUT_B620 16'hAB2E
`define CUBE_LUT_B61F 16'hAB2B
`define CUBE_LUT_B61E 16'hAB27
`define CUBE_LUT_B61D 16'hAB24
`define CUBE_LUT_B61C 16'hAB20
`define CUBE_LUT_B61B 16'hAB1D
`define CUBE_LUT_B61A 16'hAB19
`define CUBE_LUT_B619 16'hAB16
`define CUBE_LUT_B618 16'hAB12
`define CUBE_LUT_B617 16'hAB0F
`define CUBE_LUT_B616 16'hAB0B
`define CUBE_LUT_B615 16'hAB08
`define CUBE_LUT_B614 16'hAB04
`define CUBE_LUT_B613 16'hAB01
`define CUBE_LUT_B612 16'hAAFD
`define CUBE_LUT_B611 16'hAAFA
`define CUBE_LUT_B610 16'hAAF7
`define CUBE_LUT_B60F 16'hAAF3
`define CUBE_LUT_B60E 16'hAAF0
`define CUBE_LUT_B60D 16'hAAEC
`define CUBE_LUT_B60C 16'hAAE9
`define CUBE_LUT_B60B 16'hAAE5
`define CUBE_LUT_B60A 16'hAAE2
`define CUBE_LUT_B609 16'hAADF
`define CUBE_LUT_B608 16'hAADB
`define CUBE_LUT_B607 16'hAAD8
`define CUBE_LUT_B606 16'hAAD4
`define CUBE_LUT_B605 16'hAAD1
`define CUBE_LUT_B604 16'hAACE
`define CUBE_LUT_B603 16'hAACA
`define CUBE_LUT_B602 16'hAAC7
`define CUBE_LUT_B601 16'hAAC3
`define CUBE_LUT_B600 16'hAAC0
`define CUBE_LUT_B5FF 16'hAABD
`define CUBE_LUT_B5FE 16'hAAB9
`define CUBE_LUT_B5FD 16'hAAB6
`define CUBE_LUT_B5FC 16'hAAB3
`define CUBE_LUT_B5FB 16'hAAAF
`define CUBE_LUT_B5FA 16'hAAAC
`define CUBE_LUT_B5F9 16'hAAA8
`define CUBE_LUT_B5F8 16'hAAA5
`define CUBE_LUT_B5F7 16'hAAA2
`define CUBE_LUT_B5F6 16'hAA9E
`define CUBE_LUT_B5F5 16'hAA9B
`define CUBE_LUT_B5F4 16'hAA98
`define CUBE_LUT_B5F3 16'hAA94
`define CUBE_LUT_B5F2 16'hAA91
`define CUBE_LUT_B5F1 16'hAA8E
`define CUBE_LUT_B5F0 16'hAA8B
`define CUBE_LUT_B5EF 16'hAA87
`define CUBE_LUT_B5EE 16'hAA84
`define CUBE_LUT_B5ED 16'hAA81
`define CUBE_LUT_B5EC 16'hAA7D
`define CUBE_LUT_B5EB 16'hAA7A
`define CUBE_LUT_B5EA 16'hAA77
`define CUBE_LUT_B5E9 16'hAA74
`define CUBE_LUT_B5E8 16'hAA70
`define CUBE_LUT_B5E7 16'hAA6D
`define CUBE_LUT_B5E6 16'hAA6A
`define CUBE_LUT_B5E5 16'hAA66
`define CUBE_LUT_B5E4 16'hAA63
`define CUBE_LUT_B5E3 16'hAA60
`define CUBE_LUT_B5E2 16'hAA5D
`define CUBE_LUT_B5E1 16'hAA59
`define CUBE_LUT_B5E0 16'hAA56
`define CUBE_LUT_B5DF 16'hAA53
`define CUBE_LUT_B5DE 16'hAA50
`define CUBE_LUT_B5DD 16'hAA4D
`define CUBE_LUT_B5DC 16'hAA49
`define CUBE_LUT_B5DB 16'hAA46
`define CUBE_LUT_B5DA 16'hAA43
`define CUBE_LUT_B5D9 16'hAA40
`define CUBE_LUT_B5D8 16'hAA3C
`define CUBE_LUT_B5D7 16'hAA39
`define CUBE_LUT_B5D6 16'hAA36
`define CUBE_LUT_B5D5 16'hAA33
`define CUBE_LUT_B5D4 16'hAA30
`define CUBE_LUT_B5D3 16'hAA2D
`define CUBE_LUT_B5D2 16'hAA29
`define CUBE_LUT_B5D1 16'hAA26
`define CUBE_LUT_B5D0 16'hAA23
`define CUBE_LUT_B5CF 16'hAA20
`define CUBE_LUT_B5CE 16'hAA1D
`define CUBE_LUT_B5CD 16'hAA1A
`define CUBE_LUT_B5CC 16'hAA16
`define CUBE_LUT_B5CB 16'hAA13
`define CUBE_LUT_B5CA 16'hAA10
`define CUBE_LUT_B5C9 16'hAA0D
`define CUBE_LUT_B5C8 16'hAA0A
`define CUBE_LUT_B5C7 16'hAA07
`define CUBE_LUT_B5C6 16'hAA04
`define CUBE_LUT_B5C5 16'hAA00
`define CUBE_LUT_B5C4 16'hA9FD
`define CUBE_LUT_B5C3 16'hA9FA
`define CUBE_LUT_B5C2 16'hA9F7
`define CUBE_LUT_B5C1 16'hA9F4
`define CUBE_LUT_B5C0 16'hA9F1
`define CUBE_LUT_B5BF 16'hA9EE
`define CUBE_LUT_B5BE 16'hA9EB
`define CUBE_LUT_B5BD 16'hA9E8
`define CUBE_LUT_B5BC 16'hA9E5
`define CUBE_LUT_B5BB 16'hA9E1
`define CUBE_LUT_B5BA 16'hA9DE
`define CUBE_LUT_B5B9 16'hA9DB
`define CUBE_LUT_B5B8 16'hA9D8
`define CUBE_LUT_B5B7 16'hA9D5
`define CUBE_LUT_B5B6 16'hA9D2
`define CUBE_LUT_B5B5 16'hA9CF
`define CUBE_LUT_B5B4 16'hA9CC
`define CUBE_LUT_B5B3 16'hA9C9
`define CUBE_LUT_B5B2 16'hA9C6
`define CUBE_LUT_B5B1 16'hA9C3
`define CUBE_LUT_B5B0 16'hA9C0
`define CUBE_LUT_B5AF 16'hA9BD
`define CUBE_LUT_B5AE 16'hA9BA
`define CUBE_LUT_B5AD 16'hA9B7
`define CUBE_LUT_B5AC 16'hA9B4
`define CUBE_LUT_B5AB 16'hA9B1
`define CUBE_LUT_B5AA 16'hA9AE
`define CUBE_LUT_B5A9 16'hA9AB
`define CUBE_LUT_B5A8 16'hA9A8
`define CUBE_LUT_B5A7 16'hA9A5
`define CUBE_LUT_B5A6 16'hA9A2
`define CUBE_LUT_B5A5 16'hA99F
`define CUBE_LUT_B5A4 16'hA99C
`define CUBE_LUT_B5A3 16'hA999
`define CUBE_LUT_B5A2 16'hA996
`define CUBE_LUT_B5A1 16'hA993
`define CUBE_LUT_B5A0 16'hA990
`define CUBE_LUT_B59F 16'hA98D
`define CUBE_LUT_B59E 16'hA98A
`define CUBE_LUT_B59D 16'hA987
`define CUBE_LUT_B59C 16'hA984
`define CUBE_LUT_B59B 16'hA981
`define CUBE_LUT_B59A 16'hA97E
`define CUBE_LUT_B599 16'hA97B
`define CUBE_LUT_B598 16'hA978
`define CUBE_LUT_B597 16'hA975
`define CUBE_LUT_B596 16'hA972
`define CUBE_LUT_B595 16'hA96F
`define CUBE_LUT_B594 16'hA96D
`define CUBE_LUT_B593 16'hA96A
`define CUBE_LUT_B592 16'hA967
`define CUBE_LUT_B591 16'hA964
`define CUBE_LUT_B590 16'hA961
`define CUBE_LUT_B58F 16'hA95E
`define CUBE_LUT_B58E 16'hA95B
`define CUBE_LUT_B58D 16'hA958
`define CUBE_LUT_B58C 16'hA955
`define CUBE_LUT_B58B 16'hA952
`define CUBE_LUT_B58A 16'hA950
`define CUBE_LUT_B589 16'hA94D
`define CUBE_LUT_B588 16'hA94A
`define CUBE_LUT_B587 16'hA947
`define CUBE_LUT_B586 16'hA944
`define CUBE_LUT_B585 16'hA941
`define CUBE_LUT_B584 16'hA93E
`define CUBE_LUT_B583 16'hA93C
`define CUBE_LUT_B582 16'hA939
`define CUBE_LUT_B581 16'hA936
`define CUBE_LUT_B580 16'hA933
`define CUBE_LUT_B57F 16'hA930
`define CUBE_LUT_B57E 16'hA92D
`define CUBE_LUT_B57D 16'hA92B
`define CUBE_LUT_B57C 16'hA928
`define CUBE_LUT_B57B 16'hA925
`define CUBE_LUT_B57A 16'hA922
`define CUBE_LUT_B579 16'hA91F
`define CUBE_LUT_B578 16'hA91C
`define CUBE_LUT_B577 16'hA91A
`define CUBE_LUT_B576 16'hA917
`define CUBE_LUT_B575 16'hA914
`define CUBE_LUT_B574 16'hA911
`define CUBE_LUT_B573 16'hA90E
`define CUBE_LUT_B572 16'hA90C
`define CUBE_LUT_B571 16'hA909
`define CUBE_LUT_B570 16'hA906
`define CUBE_LUT_B56F 16'hA903
`define CUBE_LUT_B56E 16'hA901
`define CUBE_LUT_B56D 16'hA8FE
`define CUBE_LUT_B56C 16'hA8FB
`define CUBE_LUT_B56B 16'hA8F8
`define CUBE_LUT_B56A 16'hA8F6
`define CUBE_LUT_B569 16'hA8F3
`define CUBE_LUT_B568 16'hA8F0
`define CUBE_LUT_B567 16'hA8ED
`define CUBE_LUT_B566 16'hA8EB
`define CUBE_LUT_B565 16'hA8E8
`define CUBE_LUT_B564 16'hA8E5
`define CUBE_LUT_B563 16'hA8E2
`define CUBE_LUT_B562 16'hA8E0
`define CUBE_LUT_B561 16'hA8DD
`define CUBE_LUT_B560 16'hA8DA
`define CUBE_LUT_B55F 16'hA8D8
`define CUBE_LUT_B55E 16'hA8D5
`define CUBE_LUT_B55D 16'hA8D2
`define CUBE_LUT_B55C 16'hA8CF
`define CUBE_LUT_B55B 16'hA8CD
`define CUBE_LUT_B55A 16'hA8CA
`define CUBE_LUT_B559 16'hA8C7
`define CUBE_LUT_B558 16'hA8C5
`define CUBE_LUT_B557 16'hA8C2
`define CUBE_LUT_B556 16'hA8BF
`define CUBE_LUT_B555 16'hA8BD
`define CUBE_LUT_B554 16'hA8BA
`define CUBE_LUT_B553 16'hA8B7
`define CUBE_LUT_B552 16'hA8B5
`define CUBE_LUT_B551 16'hA8B2
`define CUBE_LUT_B550 16'hA8AF
`define CUBE_LUT_B54F 16'hA8AD
`define CUBE_LUT_B54E 16'hA8AA
`define CUBE_LUT_B54D 16'hA8A8
`define CUBE_LUT_B54C 16'hA8A5
`define CUBE_LUT_B54B 16'hA8A2
`define CUBE_LUT_B54A 16'hA8A0
`define CUBE_LUT_B549 16'hA89D
`define CUBE_LUT_B548 16'hA89A
`define CUBE_LUT_B547 16'hA898
`define CUBE_LUT_B546 16'hA895
`define CUBE_LUT_B545 16'hA893
`define CUBE_LUT_B544 16'hA890
`define CUBE_LUT_B543 16'hA88D
`define CUBE_LUT_B542 16'hA88B
`define CUBE_LUT_B541 16'hA888
`define CUBE_LUT_B540 16'hA886
`define CUBE_LUT_B53F 16'hA883
`define CUBE_LUT_B53E 16'hA880
`define CUBE_LUT_B53D 16'hA87E
`define CUBE_LUT_B53C 16'hA87B
`define CUBE_LUT_B53B 16'hA879
`define CUBE_LUT_B53A 16'hA876
`define CUBE_LUT_B539 16'hA874
`define CUBE_LUT_B538 16'hA871
`define CUBE_LUT_B537 16'hA86F
`define CUBE_LUT_B536 16'hA86C
`define CUBE_LUT_B535 16'hA869
`define CUBE_LUT_B534 16'hA867
`define CUBE_LUT_B533 16'hA864
`define CUBE_LUT_B532 16'hA862
`define CUBE_LUT_B531 16'hA85F
`define CUBE_LUT_B530 16'hA85D
`define CUBE_LUT_B52F 16'hA85A
`define CUBE_LUT_B52E 16'hA858
`define CUBE_LUT_B52D 16'hA855
`define CUBE_LUT_B52C 16'hA853
`define CUBE_LUT_B52B 16'hA850
`define CUBE_LUT_B52A 16'hA84E
`define CUBE_LUT_B529 16'hA84B
`define CUBE_LUT_B528 16'hA849
`define CUBE_LUT_B527 16'hA846
`define CUBE_LUT_B526 16'hA844
`define CUBE_LUT_B525 16'hA841
`define CUBE_LUT_B524 16'hA83F
`define CUBE_LUT_B523 16'hA83C
`define CUBE_LUT_B522 16'hA83A
`define CUBE_LUT_B521 16'hA837
`define CUBE_LUT_B520 16'hA835
`define CUBE_LUT_B51F 16'hA832
`define CUBE_LUT_B51E 16'hA830
`define CUBE_LUT_B51D 16'hA82E
`define CUBE_LUT_B51C 16'hA82B
`define CUBE_LUT_B51B 16'hA829
`define CUBE_LUT_B51A 16'hA826
`define CUBE_LUT_B519 16'hA824
`define CUBE_LUT_B518 16'hA821
`define CUBE_LUT_B517 16'hA81F
`define CUBE_LUT_B516 16'hA81C
`define CUBE_LUT_B515 16'hA81A
`define CUBE_LUT_B514 16'hA818
`define CUBE_LUT_B513 16'hA815
`define CUBE_LUT_B512 16'hA813
`define CUBE_LUT_B511 16'hA810
`define CUBE_LUT_B510 16'hA80E
`define CUBE_LUT_B50F 16'hA80C
`define CUBE_LUT_B50E 16'hA809
`define CUBE_LUT_B50D 16'hA807
`define CUBE_LUT_B50C 16'hA804
`define CUBE_LUT_B50B 16'hA802
`define CUBE_LUT_B50A 16'hA7FF
`define CUBE_LUT_B509 16'hA7FA
`define CUBE_LUT_B508 16'hA7F6
`define CUBE_LUT_B507 16'hA7F1
`define CUBE_LUT_B506 16'hA7EC
`define CUBE_LUT_B505 16'hA7E8
`define CUBE_LUT_B504 16'hA7E3
`define CUBE_LUT_B503 16'hA7DE
`define CUBE_LUT_B502 16'hA7D9
`define CUBE_LUT_B501 16'hA7D5
`define CUBE_LUT_B500 16'hA7D0
`define CUBE_LUT_B4FF 16'hA7CB
`define CUBE_LUT_B4FE 16'hA7C7
`define CUBE_LUT_B4FD 16'hA7C2
`define CUBE_LUT_B4FC 16'hA7BD
`define CUBE_LUT_B4FB 16'hA7B9
`define CUBE_LUT_B4FA 16'hA7B4
`define CUBE_LUT_B4F9 16'hA7AF
`define CUBE_LUT_B4F8 16'hA7AB
`define CUBE_LUT_B4F7 16'hA7A6
`define CUBE_LUT_B4F6 16'hA7A1
`define CUBE_LUT_B4F5 16'hA79D
`define CUBE_LUT_B4F4 16'hA798
`define CUBE_LUT_B4F3 16'hA794
`define CUBE_LUT_B4F2 16'hA78F
`define CUBE_LUT_B4F1 16'hA78B
`define CUBE_LUT_B4F0 16'hA786
`define CUBE_LUT_B4EF 16'hA781
`define CUBE_LUT_B4EE 16'hA77D
`define CUBE_LUT_B4ED 16'hA778
`define CUBE_LUT_B4EC 16'hA774
`define CUBE_LUT_B4EB 16'hA76F
`define CUBE_LUT_B4EA 16'hA76B
`define CUBE_LUT_B4E9 16'hA766
`define CUBE_LUT_B4E8 16'hA762
`define CUBE_LUT_B4E7 16'hA75D
`define CUBE_LUT_B4E6 16'hA759
`define CUBE_LUT_B4E5 16'hA754
`define CUBE_LUT_B4E4 16'hA750
`define CUBE_LUT_B4E3 16'hA74B
`define CUBE_LUT_B4E2 16'hA747
`define CUBE_LUT_B4E1 16'hA742
`define CUBE_LUT_B4E0 16'hA73E
`define CUBE_LUT_B4DF 16'hA739
`define CUBE_LUT_B4DE 16'hA735
`define CUBE_LUT_B4DD 16'hA730
`define CUBE_LUT_B4DC 16'hA72C
`define CUBE_LUT_B4DB 16'hA728
`define CUBE_LUT_B4DA 16'hA723
`define CUBE_LUT_B4D9 16'hA71F
`define CUBE_LUT_B4D8 16'hA71A
`define CUBE_LUT_B4D7 16'hA716
`define CUBE_LUT_B4D6 16'hA712
`define CUBE_LUT_B4D5 16'hA70D
`define CUBE_LUT_B4D4 16'hA709
`define CUBE_LUT_B4D3 16'hA704
`define CUBE_LUT_B4D2 16'hA700
`define CUBE_LUT_B4D1 16'hA6FC
`define CUBE_LUT_B4D0 16'hA6F7
`define CUBE_LUT_B4CF 16'hA6F3
`define CUBE_LUT_B4CE 16'hA6EF
`define CUBE_LUT_B4CD 16'hA6EA
`define CUBE_LUT_B4CC 16'hA6E6
`define CUBE_LUT_B4CB 16'hA6E2
`define CUBE_LUT_B4CA 16'hA6DD
`define CUBE_LUT_B4C9 16'hA6D9
`define CUBE_LUT_B4C8 16'hA6D5
`define CUBE_LUT_B4C7 16'hA6D1
`define CUBE_LUT_B4C6 16'hA6CC
`define CUBE_LUT_B4C5 16'hA6C8
`define CUBE_LUT_B4C4 16'hA6C4
`define CUBE_LUT_B4C3 16'hA6BF
`define CUBE_LUT_B4C2 16'hA6BB
`define CUBE_LUT_B4C1 16'hA6B7
`define CUBE_LUT_B4C0 16'hA6B3
`define CUBE_LUT_B4BF 16'hA6AF
`define CUBE_LUT_B4BE 16'hA6AA
`define CUBE_LUT_B4BD 16'hA6A6
`define CUBE_LUT_B4BC 16'hA6A2
`define CUBE_LUT_B4BB 16'hA69E
`define CUBE_LUT_B4BA 16'hA699
`define CUBE_LUT_B4B9 16'hA695
`define CUBE_LUT_B4B8 16'hA691
`define CUBE_LUT_B4B7 16'hA68D
`define CUBE_LUT_B4B6 16'hA689
`define CUBE_LUT_B4B5 16'hA685
`define CUBE_LUT_B4B4 16'hA680
`define CUBE_LUT_B4B3 16'hA67C
`define CUBE_LUT_B4B2 16'hA678
`define CUBE_LUT_B4B1 16'hA674
`define CUBE_LUT_B4B0 16'hA670
`define CUBE_LUT_B4AF 16'hA66C
`define CUBE_LUT_B4AE 16'hA668
`define CUBE_LUT_B4AD 16'hA664
`define CUBE_LUT_B4AC 16'hA660
`define CUBE_LUT_B4AB 16'hA65B
`define CUBE_LUT_B4AA 16'hA657
`define CUBE_LUT_B4A9 16'hA653
`define CUBE_LUT_B4A8 16'hA64F
`define CUBE_LUT_B4A7 16'hA64B
`define CUBE_LUT_B4A6 16'hA647
`define CUBE_LUT_B4A5 16'hA643
`define CUBE_LUT_B4A4 16'hA63F
`define CUBE_LUT_B4A3 16'hA63B
`define CUBE_LUT_B4A2 16'hA637
`define CUBE_LUT_B4A1 16'hA633
`define CUBE_LUT_B4A0 16'hA62F
`define CUBE_LUT_B49F 16'hA62B
`define CUBE_LUT_B49E 16'hA627
`define CUBE_LUT_B49D 16'hA623
`define CUBE_LUT_B49C 16'hA61F
`define CUBE_LUT_B49B 16'hA61B
`define CUBE_LUT_B49A 16'hA617
`define CUBE_LUT_B499 16'hA613
`define CUBE_LUT_B498 16'hA60F
`define CUBE_LUT_B497 16'hA60B
`define CUBE_LUT_B496 16'hA607
`define CUBE_LUT_B495 16'hA603
`define CUBE_LUT_B494 16'hA5FF
`define CUBE_LUT_B493 16'hA5FB
`define CUBE_LUT_B492 16'hA5F7
`define CUBE_LUT_B491 16'hA5F4
`define CUBE_LUT_B490 16'hA5F0
`define CUBE_LUT_B48F 16'hA5EC
`define CUBE_LUT_B48E 16'hA5E8
`define CUBE_LUT_B48D 16'hA5E4
`define CUBE_LUT_B48C 16'hA5E0
`define CUBE_LUT_B48B 16'hA5DC
`define CUBE_LUT_B48A 16'hA5D8
`define CUBE_LUT_B489 16'hA5D4
`define CUBE_LUT_B488 16'hA5D1
`define CUBE_LUT_B487 16'hA5CD
`define CUBE_LUT_B486 16'hA5C9
`define CUBE_LUT_B485 16'hA5C5
`define CUBE_LUT_B484 16'hA5C1
`define CUBE_LUT_B483 16'hA5BD
`define CUBE_LUT_B482 16'hA5BA
`define CUBE_LUT_B481 16'hA5B6
`define CUBE_LUT_B480 16'hA5B2
`define CUBE_LUT_B47F 16'hA5AE
`define CUBE_LUT_B47E 16'hA5AA
`define CUBE_LUT_B47D 16'hA5A7
`define CUBE_LUT_B47C 16'hA5A3
`define CUBE_LUT_B47B 16'hA59F
`define CUBE_LUT_B47A 16'hA59B
`define CUBE_LUT_B479 16'hA598
`define CUBE_LUT_B478 16'hA594
`define CUBE_LUT_B477 16'hA590
`define CUBE_LUT_B476 16'hA58C
`define CUBE_LUT_B475 16'hA589
`define CUBE_LUT_B474 16'hA585
`define CUBE_LUT_B473 16'hA581
`define CUBE_LUT_B472 16'hA57D
`define CUBE_LUT_B471 16'hA57A
`define CUBE_LUT_B470 16'hA576
`define CUBE_LUT_B46F 16'hA572
`define CUBE_LUT_B46E 16'hA56F
`define CUBE_LUT_B46D 16'hA56B
`define CUBE_LUT_B46C 16'hA567
`define CUBE_LUT_B46B 16'hA564
`define CUBE_LUT_B46A 16'hA560
`define CUBE_LUT_B469 16'hA55C
`define CUBE_LUT_B468 16'hA559
`define CUBE_LUT_B467 16'hA555
`define CUBE_LUT_B466 16'hA551
`define CUBE_LUT_B465 16'hA54E
`define CUBE_LUT_B464 16'hA54A
`define CUBE_LUT_B463 16'hA547
`define CUBE_LUT_B462 16'hA543
`define CUBE_LUT_B461 16'hA53F
`define CUBE_LUT_B460 16'hA53C
`define CUBE_LUT_B45F 16'hA538
`define CUBE_LUT_B45E 16'hA535
`define CUBE_LUT_B45D 16'hA531
`define CUBE_LUT_B45C 16'hA52E
`define CUBE_LUT_B45B 16'hA52A
`define CUBE_LUT_B45A 16'hA526
`define CUBE_LUT_B459 16'hA523
`define CUBE_LUT_B458 16'hA51F
`define CUBE_LUT_B457 16'hA51C
`define CUBE_LUT_B456 16'hA518
`define CUBE_LUT_B455 16'hA515
`define CUBE_LUT_B454 16'hA511
`define CUBE_LUT_B453 16'hA50E
`define CUBE_LUT_B452 16'hA50A
`define CUBE_LUT_B451 16'hA507
`define CUBE_LUT_B450 16'hA503
`define CUBE_LUT_B44F 16'hA500
`define CUBE_LUT_B44E 16'hA4FC
`define CUBE_LUT_B44D 16'hA4F9
`define CUBE_LUT_B44C 16'hA4F5
`define CUBE_LUT_B44B 16'hA4F2
`define CUBE_LUT_B44A 16'hA4EE
`define CUBE_LUT_B449 16'hA4EB
`define CUBE_LUT_B448 16'hA4E8
`define CUBE_LUT_B447 16'hA4E4
`define CUBE_LUT_B446 16'hA4E1
`define CUBE_LUT_B445 16'hA4DD
`define CUBE_LUT_B444 16'hA4DA
`define CUBE_LUT_B443 16'hA4D6
`define CUBE_LUT_B442 16'hA4D3
`define CUBE_LUT_B441 16'hA4D0
`define CUBE_LUT_B440 16'hA4CC
`define CUBE_LUT_B43F 16'hA4C9
`define CUBE_LUT_B43E 16'hA4C5
`define CUBE_LUT_B43D 16'hA4C2
`define CUBE_LUT_B43C 16'hA4BF
`define CUBE_LUT_B43B 16'hA4BB
`define CUBE_LUT_B43A 16'hA4B8
`define CUBE_LUT_B439 16'hA4B5
`define CUBE_LUT_B438 16'hA4B1
`define CUBE_LUT_B437 16'hA4AE
`define CUBE_LUT_B436 16'hA4AB
`define CUBE_LUT_B435 16'hA4A7
`define CUBE_LUT_B434 16'hA4A4
`define CUBE_LUT_B433 16'hA4A1
`define CUBE_LUT_B432 16'hA49D
`define CUBE_LUT_B431 16'hA49A
`define CUBE_LUT_B430 16'hA497
`define CUBE_LUT_B42F 16'hA494
`define CUBE_LUT_B42E 16'hA490
`define CUBE_LUT_B42D 16'hA48D
`define CUBE_LUT_B42C 16'hA48A
`define CUBE_LUT_B42B 16'hA486
`define CUBE_LUT_B42A 16'hA483
`define CUBE_LUT_B429 16'hA480
`define CUBE_LUT_B428 16'hA47D
`define CUBE_LUT_B427 16'hA47A
`define CUBE_LUT_B426 16'hA476
`define CUBE_LUT_B425 16'hA473
`define CUBE_LUT_B424 16'hA470
`define CUBE_LUT_B423 16'hA46D
`define CUBE_LUT_B422 16'hA469
`define CUBE_LUT_B421 16'hA466
`define CUBE_LUT_B420 16'hA463
`define CUBE_LUT_B41F 16'hA460
`define CUBE_LUT_B41E 16'hA45D
`define CUBE_LUT_B41D 16'hA459
`define CUBE_LUT_B41C 16'hA456
`define CUBE_LUT_B41B 16'hA453
`define CUBE_LUT_B41A 16'hA450
`define CUBE_LUT_B419 16'hA44D
`define CUBE_LUT_B418 16'hA44A
`define CUBE_LUT_B417 16'hA447
`define CUBE_LUT_B416 16'hA443
`define CUBE_LUT_B415 16'hA440
`define CUBE_LUT_B414 16'hA43D
`define CUBE_LUT_B413 16'hA43A
`define CUBE_LUT_B412 16'hA437
`define CUBE_LUT_B411 16'hA434
`define CUBE_LUT_B410 16'hA431
`define CUBE_LUT_B40F 16'hA42E
`define CUBE_LUT_B40E 16'hA42B
`define CUBE_LUT_B40D 16'hA427
`define CUBE_LUT_B40C 16'hA424
`define CUBE_LUT_B40B 16'hA421
`define CUBE_LUT_B40A 16'hA41E
`define CUBE_LUT_B409 16'hA41B
`define CUBE_LUT_B408 16'hA418
`define CUBE_LUT_B407 16'hA415
`define CUBE_LUT_B406 16'hA412
`define CUBE_LUT_B405 16'hA40F
`define CUBE_LUT_B404 16'hA40C
`define CUBE_LUT_B403 16'hA409
`define CUBE_LUT_B402 16'hA406
`define CUBE_LUT_B401 16'hA403
`define CUBE_LUT_B400 16'hA400
`define CUBE_LUT_B3FF 16'hA3FD
`define CUBE_LUT_B3FE 16'hA3FA
`define CUBE_LUT_B3FD 16'hA3F7
`define CUBE_LUT_B3FC 16'hA3F4
`define CUBE_LUT_B3FB 16'hA3F1
`define CUBE_LUT_B3FA 16'hA3EE
`define CUBE_LUT_B3F9 16'hA3EB
`define CUBE_LUT_B3F8 16'hA3E8
`define CUBE_LUT_B3F7 16'hA3E5
`define CUBE_LUT_B3F6 16'hA3E2
`define CUBE_LUT_B3F5 16'hA3DF
`define CUBE_LUT_B3F4 16'hA3DC
`define CUBE_LUT_B3F3 16'hA3D9
`define CUBE_LUT_B3F2 16'hA3D6
`define CUBE_LUT_B3F1 16'hA3D3
`define CUBE_LUT_B3F0 16'hA3D0
`define CUBE_LUT_B3EF 16'hA3CD
`define CUBE_LUT_B3EE 16'hA3CA
`define CUBE_LUT_B3ED 16'hA3C8
`define CUBE_LUT_B3EC 16'hA3C5
`define CUBE_LUT_B3EB 16'hA3C2
`define CUBE_LUT_B3EA 16'hA3BF
`define CUBE_LUT_B3E9 16'hA3BC
`define CUBE_LUT_B3E8 16'hA3B9
`define CUBE_LUT_B3E7 16'hA3B6
`define CUBE_LUT_B3E6 16'hA3B3
`define CUBE_LUT_B3E5 16'hA3B0
`define CUBE_LUT_B3E4 16'hA3AD
`define CUBE_LUT_B3E3 16'hA3AA
`define CUBE_LUT_B3E2 16'hA3A7
`define CUBE_LUT_B3E1 16'hA3A4
`define CUBE_LUT_B3E0 16'hA3A1
`define CUBE_LUT_B3DF 16'hA39F
`define CUBE_LUT_B3DE 16'hA39C
`define CUBE_LUT_B3DD 16'hA399
`define CUBE_LUT_B3DC 16'hA396
`define CUBE_LUT_B3DB 16'hA393
`define CUBE_LUT_B3DA 16'hA390
`define CUBE_LUT_B3D9 16'hA38D
`define CUBE_LUT_B3D8 16'hA38A
`define CUBE_LUT_B3D7 16'hA387
`define CUBE_LUT_B3D6 16'hA385
`define CUBE_LUT_B3D5 16'hA382
`define CUBE_LUT_B3D4 16'hA37F
`define CUBE_LUT_B3D3 16'hA37C
`define CUBE_LUT_B3D2 16'hA379
`define CUBE_LUT_B3D1 16'hA376
`define CUBE_LUT_B3D0 16'hA373
`define CUBE_LUT_B3CF 16'hA370
`define CUBE_LUT_B3CE 16'hA36E
`define CUBE_LUT_B3CD 16'hA36B
`define CUBE_LUT_B3CC 16'hA368
`define CUBE_LUT_B3CB 16'hA365
`define CUBE_LUT_B3CA 16'hA362
`define CUBE_LUT_B3C9 16'hA35F
`define CUBE_LUT_B3C8 16'hA35D
`define CUBE_LUT_B3C7 16'hA35A
`define CUBE_LUT_B3C6 16'hA357
`define CUBE_LUT_B3C5 16'hA354
`define CUBE_LUT_B3C4 16'hA351
`define CUBE_LUT_B3C3 16'hA34E
`define CUBE_LUT_B3C2 16'hA34C
`define CUBE_LUT_B3C1 16'hA349
`define CUBE_LUT_B3C0 16'hA346
`define CUBE_LUT_B3BF 16'hA343
`define CUBE_LUT_B3BE 16'hA340
`define CUBE_LUT_B3BD 16'hA33E
`define CUBE_LUT_B3BC 16'hA33B
`define CUBE_LUT_B3BB 16'hA338
`define CUBE_LUT_B3BA 16'hA335
`define CUBE_LUT_B3B9 16'hA332
`define CUBE_LUT_B3B8 16'hA330
`define CUBE_LUT_B3B7 16'hA32D
`define CUBE_LUT_B3B6 16'hA32A
`define CUBE_LUT_B3B5 16'hA327
`define CUBE_LUT_B3B4 16'hA324
`define CUBE_LUT_B3B3 16'hA322
`define CUBE_LUT_B3B2 16'hA31F
`define CUBE_LUT_B3B1 16'hA31C
`define CUBE_LUT_B3B0 16'hA319
`define CUBE_LUT_B3AF 16'hA316
`define CUBE_LUT_B3AE 16'hA314
`define CUBE_LUT_B3AD 16'hA311
`define CUBE_LUT_B3AC 16'hA30E
`define CUBE_LUT_B3AB 16'hA30B
`define CUBE_LUT_B3AA 16'hA309
`define CUBE_LUT_B3A9 16'hA306
`define CUBE_LUT_B3A8 16'hA303
`define CUBE_LUT_B3A7 16'hA300
`define CUBE_LUT_B3A6 16'hA2FE
`define CUBE_LUT_B3A5 16'hA2FB
`define CUBE_LUT_B3A4 16'hA2F8
`define CUBE_LUT_B3A3 16'hA2F5
`define CUBE_LUT_B3A2 16'hA2F3
`define CUBE_LUT_B3A1 16'hA2F0
`define CUBE_LUT_B3A0 16'hA2ED
`define CUBE_LUT_B39F 16'hA2EB
`define CUBE_LUT_B39E 16'hA2E8
`define CUBE_LUT_B39D 16'hA2E5
`define CUBE_LUT_B39C 16'hA2E2
`define CUBE_LUT_B39B 16'hA2E0
`define CUBE_LUT_B39A 16'hA2DD
`define CUBE_LUT_B399 16'hA2DA
`define CUBE_LUT_B398 16'hA2D8
`define CUBE_LUT_B397 16'hA2D5
`define CUBE_LUT_B396 16'hA2D2
`define CUBE_LUT_B395 16'hA2CF
`define CUBE_LUT_B394 16'hA2CD
`define CUBE_LUT_B393 16'hA2CA
`define CUBE_LUT_B392 16'hA2C7
`define CUBE_LUT_B391 16'hA2C5
`define CUBE_LUT_B390 16'hA2C2
`define CUBE_LUT_B38F 16'hA2BF
`define CUBE_LUT_B38E 16'hA2BD
`define CUBE_LUT_B38D 16'hA2BA
`define CUBE_LUT_B38C 16'hA2B7
`define CUBE_LUT_B38B 16'hA2B5
`define CUBE_LUT_B38A 16'hA2B2
`define CUBE_LUT_B389 16'hA2AF
`define CUBE_LUT_B388 16'hA2AD
`define CUBE_LUT_B387 16'hA2AA
`define CUBE_LUT_B386 16'hA2A7
`define CUBE_LUT_B385 16'hA2A5
`define CUBE_LUT_B384 16'hA2A2
`define CUBE_LUT_B383 16'hA29F
`define CUBE_LUT_B382 16'hA29D
`define CUBE_LUT_B381 16'hA29A
`define CUBE_LUT_B380 16'hA298
`define CUBE_LUT_B37F 16'hA295
`define CUBE_LUT_B37E 16'hA292
`define CUBE_LUT_B37D 16'hA290
`define CUBE_LUT_B37C 16'hA28D
`define CUBE_LUT_B37B 16'hA28A
`define CUBE_LUT_B37A 16'hA288
`define CUBE_LUT_B379 16'hA285
`define CUBE_LUT_B378 16'hA282
`define CUBE_LUT_B377 16'hA280
`define CUBE_LUT_B376 16'hA27D
`define CUBE_LUT_B375 16'hA27B
`define CUBE_LUT_B374 16'hA278
`define CUBE_LUT_B373 16'hA275
`define CUBE_LUT_B372 16'hA273
`define CUBE_LUT_B371 16'hA270
`define CUBE_LUT_B370 16'hA26E
`define CUBE_LUT_B36F 16'hA26B
`define CUBE_LUT_B36E 16'hA268
`define CUBE_LUT_B36D 16'hA266
`define CUBE_LUT_B36C 16'hA263
`define CUBE_LUT_B36B 16'hA261
`define CUBE_LUT_B36A 16'hA25E
`define CUBE_LUT_B369 16'hA25C
`define CUBE_LUT_B368 16'hA259
`define CUBE_LUT_B367 16'hA256
`define CUBE_LUT_B366 16'hA254
`define CUBE_LUT_B365 16'hA251
`define CUBE_LUT_B364 16'hA24F
`define CUBE_LUT_B363 16'hA24C
`define CUBE_LUT_B362 16'hA24A
`define CUBE_LUT_B361 16'hA247
`define CUBE_LUT_B360 16'hA245
`define CUBE_LUT_B35F 16'hA242
`define CUBE_LUT_B35E 16'hA23F
`define CUBE_LUT_B35D 16'hA23D
`define CUBE_LUT_B35C 16'hA23A
`define CUBE_LUT_B35B 16'hA238
`define CUBE_LUT_B35A 16'hA235
`define CUBE_LUT_B359 16'hA233
`define CUBE_LUT_B358 16'hA230
`define CUBE_LUT_B357 16'hA22E
`define CUBE_LUT_B356 16'hA22B
`define CUBE_LUT_B355 16'hA229
`define CUBE_LUT_B354 16'hA226
`define CUBE_LUT_B353 16'hA224
`define CUBE_LUT_B352 16'hA221
`define CUBE_LUT_B351 16'hA21F
`define CUBE_LUT_B350 16'hA21C
`define CUBE_LUT_B34F 16'hA21A
`define CUBE_LUT_B34E 16'hA217
`define CUBE_LUT_B34D 16'hA215
`define CUBE_LUT_B34C 16'hA212
`define CUBE_LUT_B34B 16'hA210
`define CUBE_LUT_B34A 16'hA20D
`define CUBE_LUT_B349 16'hA20B
`define CUBE_LUT_B348 16'hA208
`define CUBE_LUT_B347 16'hA206
`define CUBE_LUT_B346 16'hA203
`define CUBE_LUT_B345 16'hA201
`define CUBE_LUT_B344 16'hA1FE
`define CUBE_LUT_B343 16'hA1FC
`define CUBE_LUT_B342 16'hA1F9
`define CUBE_LUT_B341 16'hA1F7
`define CUBE_LUT_B340 16'hA1F4
`define CUBE_LUT_B33F 16'hA1F2
`define CUBE_LUT_B33E 16'hA1EF
`define CUBE_LUT_B33D 16'hA1ED
`define CUBE_LUT_B33C 16'hA1EA
`define CUBE_LUT_B33B 16'hA1E8
`define CUBE_LUT_B33A 16'hA1E6
`define CUBE_LUT_B339 16'hA1E3
`define CUBE_LUT_B338 16'hA1E1
`define CUBE_LUT_B337 16'hA1DE
`define CUBE_LUT_B336 16'hA1DC
`define CUBE_LUT_B335 16'hA1D9
`define CUBE_LUT_B334 16'hA1D7
`define CUBE_LUT_B333 16'hA1D5
`define CUBE_LUT_B332 16'hA1D2
`define CUBE_LUT_B331 16'hA1D0
`define CUBE_LUT_B330 16'hA1CD
`define CUBE_LUT_B32F 16'hA1CB
`define CUBE_LUT_B32E 16'hA1C8
`define CUBE_LUT_B32D 16'hA1C6
`define CUBE_LUT_B32C 16'hA1C4
`define CUBE_LUT_B32B 16'hA1C1
`define CUBE_LUT_B32A 16'hA1BF
`define CUBE_LUT_B329 16'hA1BC
`define CUBE_LUT_B328 16'hA1BA
`define CUBE_LUT_B327 16'hA1B8
`define CUBE_LUT_B326 16'hA1B5
`define CUBE_LUT_B325 16'hA1B3
`define CUBE_LUT_B324 16'hA1B0
`define CUBE_LUT_B323 16'hA1AE
`define CUBE_LUT_B322 16'hA1AC
`define CUBE_LUT_B321 16'hA1A9
`define CUBE_LUT_B320 16'hA1A7
`define CUBE_LUT_B31F 16'hA1A4
`define CUBE_LUT_B31E 16'hA1A2
`define CUBE_LUT_B31D 16'hA1A0
`define CUBE_LUT_B31C 16'hA19D
`define CUBE_LUT_B31B 16'hA19B
`define CUBE_LUT_B31A 16'hA199
`define CUBE_LUT_B319 16'hA196
`define CUBE_LUT_B318 16'hA194
`define CUBE_LUT_B317 16'hA192
`define CUBE_LUT_B316 16'hA18F
`define CUBE_LUT_B315 16'hA18D
`define CUBE_LUT_B314 16'hA18A
`define CUBE_LUT_B313 16'hA188
`define CUBE_LUT_B312 16'hA186
`define CUBE_LUT_B311 16'hA183
`define CUBE_LUT_B310 16'hA181
`define CUBE_LUT_B30F 16'hA17F
`define CUBE_LUT_B30E 16'hA17C
`define CUBE_LUT_B30D 16'hA17A
`define CUBE_LUT_B30C 16'hA178
`define CUBE_LUT_B30B 16'hA175
`define CUBE_LUT_B30A 16'hA173
`define CUBE_LUT_B309 16'hA171
`define CUBE_LUT_B308 16'hA16E
`define CUBE_LUT_B307 16'hA16C
`define CUBE_LUT_B306 16'hA16A
`define CUBE_LUT_B305 16'hA168
`define CUBE_LUT_B304 16'hA165
`define CUBE_LUT_B303 16'hA163
`define CUBE_LUT_B302 16'hA161
`define CUBE_LUT_B301 16'hA15E
`define CUBE_LUT_B300 16'hA15C
`define CUBE_LUT_B2FF 16'hA15A
`define CUBE_LUT_B2FE 16'hA157
`define CUBE_LUT_B2FD 16'hA155
`define CUBE_LUT_B2FC 16'hA153
`define CUBE_LUT_B2FB 16'hA151
`define CUBE_LUT_B2FA 16'hA14E
`define CUBE_LUT_B2F9 16'hA14C
`define CUBE_LUT_B2F8 16'hA14A
`define CUBE_LUT_B2F7 16'hA147
`define CUBE_LUT_B2F6 16'hA145
`define CUBE_LUT_B2F5 16'hA143
`define CUBE_LUT_B2F4 16'hA141
`define CUBE_LUT_B2F3 16'hA13E
`define CUBE_LUT_B2F2 16'hA13C
`define CUBE_LUT_B2F1 16'hA13A
`define CUBE_LUT_B2F0 16'hA138
`define CUBE_LUT_B2EF 16'hA135
`define CUBE_LUT_B2EE 16'hA133
`define CUBE_LUT_B2ED 16'hA131
`define CUBE_LUT_B2EC 16'hA12F
`define CUBE_LUT_B2EB 16'hA12C
`define CUBE_LUT_B2EA 16'hA12A
`define CUBE_LUT_B2E9 16'hA128
`define CUBE_LUT_B2E8 16'hA126
`define CUBE_LUT_B2E7 16'hA123
`define CUBE_LUT_B2E6 16'hA121
`define CUBE_LUT_B2E5 16'hA11F
`define CUBE_LUT_B2E4 16'hA11D
`define CUBE_LUT_B2E3 16'hA11A
`define CUBE_LUT_B2E2 16'hA118
`define CUBE_LUT_B2E1 16'hA116
`define CUBE_LUT_B2E0 16'hA114
`define CUBE_LUT_B2DF 16'hA112
`define CUBE_LUT_B2DE 16'hA10F
`define CUBE_LUT_B2DD 16'hA10D
`define CUBE_LUT_B2DC 16'hA10B
`define CUBE_LUT_B2DB 16'hA109
`define CUBE_LUT_B2DA 16'hA107
`define CUBE_LUT_B2D9 16'hA104
`define CUBE_LUT_B2D8 16'hA102
`define CUBE_LUT_B2D7 16'hA100
`define CUBE_LUT_B2D6 16'hA0FE
`define CUBE_LUT_B2D5 16'hA0FC
`define CUBE_LUT_B2D4 16'hA0F9
`define CUBE_LUT_B2D3 16'hA0F7
`define CUBE_LUT_B2D2 16'hA0F5
`define CUBE_LUT_B2D1 16'hA0F3
`define CUBE_LUT_B2D0 16'hA0F1
`define CUBE_LUT_B2CF 16'hA0EF
`define CUBE_LUT_B2CE 16'hA0EC
`define CUBE_LUT_B2CD 16'hA0EA
`define CUBE_LUT_B2CC 16'hA0E8
`define CUBE_LUT_B2CB 16'hA0E6
`define CUBE_LUT_B2CA 16'hA0E4
`define CUBE_LUT_B2C9 16'hA0E2
`define CUBE_LUT_B2C8 16'hA0DF
`define CUBE_LUT_B2C7 16'hA0DD
`define CUBE_LUT_B2C6 16'hA0DB
`define CUBE_LUT_B2C5 16'hA0D9
`define CUBE_LUT_B2C4 16'hA0D7
`define CUBE_LUT_B2C3 16'hA0D5
`define CUBE_LUT_B2C2 16'hA0D2
`define CUBE_LUT_B2C1 16'hA0D0
`define CUBE_LUT_B2C0 16'hA0CE
`define CUBE_LUT_B2BF 16'hA0CC
`define CUBE_LUT_B2BE 16'hA0CA
`define CUBE_LUT_B2BD 16'hA0C8
`define CUBE_LUT_B2BC 16'hA0C6
`define CUBE_LUT_B2BB 16'hA0C4
`define CUBE_LUT_B2BA 16'hA0C1
`define CUBE_LUT_B2B9 16'hA0BF
`define CUBE_LUT_B2B8 16'hA0BD
`define CUBE_LUT_B2B7 16'hA0BB
`define CUBE_LUT_B2B6 16'hA0B9
`define CUBE_LUT_B2B5 16'hA0B7
`define CUBE_LUT_B2B4 16'hA0B5
`define CUBE_LUT_B2B3 16'hA0B3
`define CUBE_LUT_B2B2 16'hA0B1
`define CUBE_LUT_B2B1 16'hA0AE
`define CUBE_LUT_B2B0 16'hA0AC
`define CUBE_LUT_B2AF 16'hA0AA
`define CUBE_LUT_B2AE 16'hA0A8
`define CUBE_LUT_B2AD 16'hA0A6
`define CUBE_LUT_B2AC 16'hA0A4
`define CUBE_LUT_B2AB 16'hA0A2
`define CUBE_LUT_B2AA 16'hA0A0
`define CUBE_LUT_B2A9 16'hA09E
`define CUBE_LUT_B2A8 16'hA09C
`define CUBE_LUT_B2A7 16'hA09A
`define CUBE_LUT_B2A6 16'hA097
`define CUBE_LUT_B2A5 16'hA095
`define CUBE_LUT_B2A4 16'hA093
`define CUBE_LUT_B2A3 16'hA091
`define CUBE_LUT_B2A2 16'hA08F
`define CUBE_LUT_B2A1 16'hA08D
`define CUBE_LUT_B2A0 16'hA08B
`define CUBE_LUT_B29F 16'hA089
`define CUBE_LUT_B29E 16'hA087
`define CUBE_LUT_B29D 16'hA085
`define CUBE_LUT_B29C 16'hA083
`define CUBE_LUT_B29B 16'hA081
`define CUBE_LUT_B29A 16'hA07F
`define CUBE_LUT_B299 16'hA07D
`define CUBE_LUT_B298 16'hA07B
`define CUBE_LUT_B297 16'hA079
`define CUBE_LUT_B296 16'hA077
`define CUBE_LUT_B295 16'hA075
`define CUBE_LUT_B294 16'hA073
`define CUBE_LUT_B293 16'hA071
`define CUBE_LUT_B292 16'hA06F
`define CUBE_LUT_B291 16'hA06D
`define CUBE_LUT_B290 16'hA06A
`define CUBE_LUT_B28F 16'hA068
`define CUBE_LUT_B28E 16'hA066
`define CUBE_LUT_B28D 16'hA064
`define CUBE_LUT_B28C 16'hA062
`define CUBE_LUT_B28B 16'hA060
`define CUBE_LUT_B28A 16'hA05E
`define CUBE_LUT_B289 16'hA05C
`define CUBE_LUT_B288 16'hA05A
`define CUBE_LUT_B287 16'hA058
`define CUBE_LUT_B286 16'hA056
`define CUBE_LUT_B285 16'hA054
`define CUBE_LUT_B284 16'hA052
`define CUBE_LUT_B283 16'hA050
`define CUBE_LUT_B282 16'hA04E
`define CUBE_LUT_B281 16'hA04C
`define CUBE_LUT_B280 16'hA04A
`define CUBE_LUT_B27F 16'hA049
`define CUBE_LUT_B27E 16'hA047
`define CUBE_LUT_B27D 16'hA045
`define CUBE_LUT_B27C 16'hA043
`define CUBE_LUT_B27B 16'hA041
`define CUBE_LUT_B27A 16'hA03F
`define CUBE_LUT_B279 16'hA03D
`define CUBE_LUT_B278 16'hA03B
`define CUBE_LUT_B277 16'hA039
`define CUBE_LUT_B276 16'hA037
`define CUBE_LUT_B275 16'hA035
`define CUBE_LUT_B274 16'hA033
`define CUBE_LUT_B273 16'hA031
`define CUBE_LUT_B272 16'hA02F
`define CUBE_LUT_B271 16'hA02D
`define CUBE_LUT_B270 16'hA02B
`define CUBE_LUT_B26F 16'hA029
`define CUBE_LUT_B26E 16'hA027
`define CUBE_LUT_B26D 16'hA025
`define CUBE_LUT_B26C 16'hA023
`define CUBE_LUT_B26B 16'hA021
`define CUBE_LUT_B26A 16'hA020
`define CUBE_LUT_B269 16'hA01E
`define CUBE_LUT_B268 16'hA01C
`define CUBE_LUT_B267 16'hA01A
`define CUBE_LUT_B266 16'hA018
`define CUBE_LUT_B265 16'hA016
`define CUBE_LUT_B264 16'hA014
`define CUBE_LUT_B263 16'hA012
`define CUBE_LUT_B262 16'hA010
`define CUBE_LUT_B261 16'hA00E
`define CUBE_LUT_B260 16'hA00C
`define CUBE_LUT_B25F 16'hA00A
`define CUBE_LUT_B25E 16'hA009
`define CUBE_LUT_B25D 16'hA007
`define CUBE_LUT_B25C 16'hA005
`define CUBE_LUT_B25B 16'hA003
`define CUBE_LUT_B25A 16'hA001
`define CUBE_LUT_B259 16'h9FFE
`define CUBE_LUT_B258 16'h9FFA
`define CUBE_LUT_B257 16'h9FF7
`define CUBE_LUT_B256 16'h9FF3
`define CUBE_LUT_B255 16'h9FEF
`define CUBE_LUT_B254 16'h9FEB
`define CUBE_LUT_B253 16'h9FE8
`define CUBE_LUT_B252 16'h9FE4
`define CUBE_LUT_B251 16'h9FE0
`define CUBE_LUT_B250 16'h9FDC
`define CUBE_LUT_B24F 16'h9FD9
`define CUBE_LUT_B24E 16'h9FD5
`define CUBE_LUT_B24D 16'h9FD1
`define CUBE_LUT_B24C 16'h9FCD
`define CUBE_LUT_B24B 16'h9FCA
`define CUBE_LUT_B24A 16'h9FC6
`define CUBE_LUT_B249 16'h9FC2
`define CUBE_LUT_B248 16'h9FBF
`define CUBE_LUT_B247 16'h9FBB
`define CUBE_LUT_B246 16'h9FB7
`define CUBE_LUT_B245 16'h9FB3
`define CUBE_LUT_B244 16'h9FB0
`define CUBE_LUT_B243 16'h9FAC
`define CUBE_LUT_B242 16'h9FA8
`define CUBE_LUT_B241 16'h9FA5
`define CUBE_LUT_B240 16'h9FA1
`define CUBE_LUT_B23F 16'h9F9D
`define CUBE_LUT_B23E 16'h9F9A
`define CUBE_LUT_B23D 16'h9F96
`define CUBE_LUT_B23C 16'h9F93
`define CUBE_LUT_B23B 16'h9F8F
`define CUBE_LUT_B23A 16'h9F8B
`define CUBE_LUT_B239 16'h9F88
`define CUBE_LUT_B238 16'h9F84
`define CUBE_LUT_B237 16'h9F80
`define CUBE_LUT_B236 16'h9F7D
`define CUBE_LUT_B235 16'h9F79
`define CUBE_LUT_B234 16'h9F76
`define CUBE_LUT_B233 16'h9F72
`define CUBE_LUT_B232 16'h9F6E
`define CUBE_LUT_B231 16'h9F6B
`define CUBE_LUT_B230 16'h9F67
`define CUBE_LUT_B22F 16'h9F64
`define CUBE_LUT_B22E 16'h9F60
`define CUBE_LUT_B22D 16'h9F5C
`define CUBE_LUT_B22C 16'h9F59
`define CUBE_LUT_B22B 16'h9F55
`define CUBE_LUT_B22A 16'h9F52
`define CUBE_LUT_B229 16'h9F4E
`define CUBE_LUT_B228 16'h9F4B
`define CUBE_LUT_B227 16'h9F47
`define CUBE_LUT_B226 16'h9F43
`define CUBE_LUT_B225 16'h9F40
`define CUBE_LUT_B224 16'h9F3C
`define CUBE_LUT_B223 16'h9F39
`define CUBE_LUT_B222 16'h9F35
`define CUBE_LUT_B221 16'h9F32
`define CUBE_LUT_B220 16'h9F2E
`define CUBE_LUT_B21F 16'h9F2B
`define CUBE_LUT_B21E 16'h9F27
`define CUBE_LUT_B21D 16'h9F24
`define CUBE_LUT_B21C 16'h9F20
`define CUBE_LUT_B21B 16'h9F1D
`define CUBE_LUT_B21A 16'h9F19
`define CUBE_LUT_B219 16'h9F16
`define CUBE_LUT_B218 16'h9F12
`define CUBE_LUT_B217 16'h9F0F
`define CUBE_LUT_B216 16'h9F0B
`define CUBE_LUT_B215 16'h9F08
`define CUBE_LUT_B214 16'h9F04
`define CUBE_LUT_B213 16'h9F01
`define CUBE_LUT_B212 16'h9EFD
`define CUBE_LUT_B211 16'h9EFA
`define CUBE_LUT_B210 16'h9EF7
`define CUBE_LUT_B20F 16'h9EF3
`define CUBE_LUT_B20E 16'h9EF0
`define CUBE_LUT_B20D 16'h9EEC
`define CUBE_LUT_B20C 16'h9EE9
`define CUBE_LUT_B20B 16'h9EE5
`define CUBE_LUT_B20A 16'h9EE2
`define CUBE_LUT_B209 16'h9EDF
`define CUBE_LUT_B208 16'h9EDB
`define CUBE_LUT_B207 16'h9ED8
`define CUBE_LUT_B206 16'h9ED4
`define CUBE_LUT_B205 16'h9ED1
`define CUBE_LUT_B204 16'h9ECE
`define CUBE_LUT_B203 16'h9ECA
`define CUBE_LUT_B202 16'h9EC7
`define CUBE_LUT_B201 16'h9EC3
`define CUBE_LUT_B200 16'h9EC0
`define CUBE_LUT_B1FF 16'h9EBD
`define CUBE_LUT_B1FE 16'h9EB9
`define CUBE_LUT_B1FD 16'h9EB6
`define CUBE_LUT_B1FC 16'h9EB3
`define CUBE_LUT_B1FB 16'h9EAF
`define CUBE_LUT_B1FA 16'h9EAC
`define CUBE_LUT_B1F9 16'h9EA8
`define CUBE_LUT_B1F8 16'h9EA5
`define CUBE_LUT_B1F7 16'h9EA2
`define CUBE_LUT_B1F6 16'h9E9E
`define CUBE_LUT_B1F5 16'h9E9B
`define CUBE_LUT_B1F4 16'h9E98
`define CUBE_LUT_B1F3 16'h9E94
`define CUBE_LUT_B1F2 16'h9E91
`define CUBE_LUT_B1F1 16'h9E8E
`define CUBE_LUT_B1F0 16'h9E8B
`define CUBE_LUT_B1EF 16'h9E87
`define CUBE_LUT_B1EE 16'h9E84
`define CUBE_LUT_B1ED 16'h9E81
`define CUBE_LUT_B1EC 16'h9E7D
`define CUBE_LUT_B1EB 16'h9E7A
`define CUBE_LUT_B1EA 16'h9E77
`define CUBE_LUT_B1E9 16'h9E74
`define CUBE_LUT_B1E8 16'h9E70
`define CUBE_LUT_B1E7 16'h9E6D
`define CUBE_LUT_B1E6 16'h9E6A
`define CUBE_LUT_B1E5 16'h9E66
`define CUBE_LUT_B1E4 16'h9E63
`define CUBE_LUT_B1E3 16'h9E60
`define CUBE_LUT_B1E2 16'h9E5D
`define CUBE_LUT_B1E1 16'h9E59
`define CUBE_LUT_B1E0 16'h9E56
`define CUBE_LUT_B1DF 16'h9E53
`define CUBE_LUT_B1DE 16'h9E50
`define CUBE_LUT_B1DD 16'h9E4D
`define CUBE_LUT_B1DC 16'h9E49
`define CUBE_LUT_B1DB 16'h9E46
`define CUBE_LUT_B1DA 16'h9E43
`define CUBE_LUT_B1D9 16'h9E40
`define CUBE_LUT_B1D8 16'h9E3C
`define CUBE_LUT_B1D7 16'h9E39
`define CUBE_LUT_B1D6 16'h9E36
`define CUBE_LUT_B1D5 16'h9E33
`define CUBE_LUT_B1D4 16'h9E30
`define CUBE_LUT_B1D3 16'h9E2D
`define CUBE_LUT_B1D2 16'h9E29
`define CUBE_LUT_B1D1 16'h9E26
`define CUBE_LUT_B1D0 16'h9E23
`define CUBE_LUT_B1CF 16'h9E20
`define CUBE_LUT_B1CE 16'h9E1D
`define CUBE_LUT_B1CD 16'h9E1A
`define CUBE_LUT_B1CC 16'h9E16
`define CUBE_LUT_B1CB 16'h9E13
`define CUBE_LUT_B1CA 16'h9E10
`define CUBE_LUT_B1C9 16'h9E0D
`define CUBE_LUT_B1C8 16'h9E0A
`define CUBE_LUT_B1C7 16'h9E07
`define CUBE_LUT_B1C6 16'h9E04
`define CUBE_LUT_B1C5 16'h9E00
`define CUBE_LUT_B1C4 16'h9DFD
`define CUBE_LUT_B1C3 16'h9DFA
`define CUBE_LUT_B1C2 16'h9DF7
`define CUBE_LUT_B1C1 16'h9DF4
`define CUBE_LUT_B1C0 16'h9DF1
`define CUBE_LUT_B1BF 16'h9DEE
`define CUBE_LUT_B1BE 16'h9DEB
`define CUBE_LUT_B1BD 16'h9DE8
`define CUBE_LUT_B1BC 16'h9DE5
`define CUBE_LUT_B1BB 16'h9DE1
`define CUBE_LUT_B1BA 16'h9DDE
`define CUBE_LUT_B1B9 16'h9DDB
`define CUBE_LUT_B1B8 16'h9DD8
`define CUBE_LUT_B1B7 16'h9DD5
`define CUBE_LUT_B1B6 16'h9DD2
`define CUBE_LUT_B1B5 16'h9DCF
`define CUBE_LUT_B1B4 16'h9DCC
`define CUBE_LUT_B1B3 16'h9DC9
`define CUBE_LUT_B1B2 16'h9DC6
`define CUBE_LUT_B1B1 16'h9DC3
`define CUBE_LUT_B1B0 16'h9DC0
`define CUBE_LUT_B1AF 16'h9DBD
`define CUBE_LUT_B1AE 16'h9DBA
`define CUBE_LUT_B1AD 16'h9DB7
`define CUBE_LUT_B1AC 16'h9DB4
`define CUBE_LUT_B1AB 16'h9DB1
`define CUBE_LUT_B1AA 16'h9DAE
`define CUBE_LUT_B1A9 16'h9DAB
`define CUBE_LUT_B1A8 16'h9DA8
`define CUBE_LUT_B1A7 16'h9DA5
`define CUBE_LUT_B1A6 16'h9DA2
`define CUBE_LUT_B1A5 16'h9D9F
`define CUBE_LUT_B1A4 16'h9D9C
`define CUBE_LUT_B1A3 16'h9D99
`define CUBE_LUT_B1A2 16'h9D96
`define CUBE_LUT_B1A1 16'h9D93
`define CUBE_LUT_B1A0 16'h9D90
`define CUBE_LUT_B19F 16'h9D8D
`define CUBE_LUT_B19E 16'h9D8A
`define CUBE_LUT_B19D 16'h9D87
`define CUBE_LUT_B19C 16'h9D84
`define CUBE_LUT_B19B 16'h9D81
`define CUBE_LUT_B19A 16'h9D7E
`define CUBE_LUT_B199 16'h9D7B
`define CUBE_LUT_B198 16'h9D78
`define CUBE_LUT_B197 16'h9D75
`define CUBE_LUT_B196 16'h9D72
`define CUBE_LUT_B195 16'h9D6F
`define CUBE_LUT_B194 16'h9D6D
`define CUBE_LUT_B193 16'h9D6A
`define CUBE_LUT_B192 16'h9D67
`define CUBE_LUT_B191 16'h9D64
`define CUBE_LUT_B190 16'h9D61
`define CUBE_LUT_B18F 16'h9D5E
`define CUBE_LUT_B18E 16'h9D5B
`define CUBE_LUT_B18D 16'h9D58
`define CUBE_LUT_B18C 16'h9D55
`define CUBE_LUT_B18B 16'h9D52
`define CUBE_LUT_B18A 16'h9D50
`define CUBE_LUT_B189 16'h9D4D
`define CUBE_LUT_B188 16'h9D4A
`define CUBE_LUT_B187 16'h9D47
`define CUBE_LUT_B186 16'h9D44
`define CUBE_LUT_B185 16'h9D41
`define CUBE_LUT_B184 16'h9D3E
`define CUBE_LUT_B183 16'h9D3C
`define CUBE_LUT_B182 16'h9D39
`define CUBE_LUT_B181 16'h9D36
`define CUBE_LUT_B180 16'h9D33
`define CUBE_LUT_B17F 16'h9D30
`define CUBE_LUT_B17E 16'h9D2D
`define CUBE_LUT_B17D 16'h9D2B
`define CUBE_LUT_B17C 16'h9D28
`define CUBE_LUT_B17B 16'h9D25
`define CUBE_LUT_B17A 16'h9D22
`define CUBE_LUT_B179 16'h9D1F
`define CUBE_LUT_B178 16'h9D1C
`define CUBE_LUT_B177 16'h9D1A
`define CUBE_LUT_B176 16'h9D17
`define CUBE_LUT_B175 16'h9D14
`define CUBE_LUT_B174 16'h9D11
`define CUBE_LUT_B173 16'h9D0E
`define CUBE_LUT_B172 16'h9D0C
`define CUBE_LUT_B171 16'h9D09
`define CUBE_LUT_B170 16'h9D06
`define CUBE_LUT_B16F 16'h9D03
`define CUBE_LUT_B16E 16'h9D01
`define CUBE_LUT_B16D 16'h9CFE
`define CUBE_LUT_B16C 16'h9CFB
`define CUBE_LUT_B16B 16'h9CF8
`define CUBE_LUT_B16A 16'h9CF6
`define CUBE_LUT_B169 16'h9CF3
`define CUBE_LUT_B168 16'h9CF0
`define CUBE_LUT_B167 16'h9CED
`define CUBE_LUT_B166 16'h9CEB
`define CUBE_LUT_B165 16'h9CE8
`define CUBE_LUT_B164 16'h9CE5
`define CUBE_LUT_B163 16'h9CE2
`define CUBE_LUT_B162 16'h9CE0
`define CUBE_LUT_B161 16'h9CDD
`define CUBE_LUT_B160 16'h9CDA
`define CUBE_LUT_B15F 16'h9CD8
`define CUBE_LUT_B15E 16'h9CD5
`define CUBE_LUT_B15D 16'h9CD2
`define CUBE_LUT_B15C 16'h9CCF
`define CUBE_LUT_B15B 16'h9CCD
`define CUBE_LUT_B15A 16'h9CCA
`define CUBE_LUT_B159 16'h9CC7
`define CUBE_LUT_B158 16'h9CC5
`define CUBE_LUT_B157 16'h9CC2
`define CUBE_LUT_B156 16'h9CBF
`define CUBE_LUT_B155 16'h9CBD
`define CUBE_LUT_B154 16'h9CBA
`define CUBE_LUT_B153 16'h9CB7
`define CUBE_LUT_B152 16'h9CB5
`define CUBE_LUT_B151 16'h9CB2
`define CUBE_LUT_B150 16'h9CAF
`define CUBE_LUT_B14F 16'h9CAD
`define CUBE_LUT_B14E 16'h9CAA
`define CUBE_LUT_B14D 16'h9CA8
`define CUBE_LUT_B14C 16'h9CA5
`define CUBE_LUT_B14B 16'h9CA2
`define CUBE_LUT_B14A 16'h9CA0
`define CUBE_LUT_B149 16'h9C9D
`define CUBE_LUT_B148 16'h9C9A
`define CUBE_LUT_B147 16'h9C98
`define CUBE_LUT_B146 16'h9C95
`define CUBE_LUT_B145 16'h9C93
`define CUBE_LUT_B144 16'h9C90
`define CUBE_LUT_B143 16'h9C8D
`define CUBE_LUT_B142 16'h9C8B
`define CUBE_LUT_B141 16'h9C88
`define CUBE_LUT_B140 16'h9C86
`define CUBE_LUT_B13F 16'h9C83
`define CUBE_LUT_B13E 16'h9C80
`define CUBE_LUT_B13D 16'h9C7E
`define CUBE_LUT_B13C 16'h9C7B
`define CUBE_LUT_B13B 16'h9C79
`define CUBE_LUT_B13A 16'h9C76
`define CUBE_LUT_B139 16'h9C74
`define CUBE_LUT_B138 16'h9C71
`define CUBE_LUT_B137 16'h9C6F
`define CUBE_LUT_B136 16'h9C6C
`define CUBE_LUT_B135 16'h9C69
`define CUBE_LUT_B134 16'h9C67
`define CUBE_LUT_B133 16'h9C64
`define CUBE_LUT_B132 16'h9C62
`define CUBE_LUT_B131 16'h9C5F
`define CUBE_LUT_B130 16'h9C5D
`define CUBE_LUT_B12F 16'h9C5A
`define CUBE_LUT_B12E 16'h9C58
`define CUBE_LUT_B12D 16'h9C55
`define CUBE_LUT_B12C 16'h9C53
`define CUBE_LUT_B12B 16'h9C50
`define CUBE_LUT_B12A 16'h9C4E
`define CUBE_LUT_B129 16'h9C4B
`define CUBE_LUT_B128 16'h9C49
`define CUBE_LUT_B127 16'h9C46
`define CUBE_LUT_B126 16'h9C44
`define CUBE_LUT_B125 16'h9C41
`define CUBE_LUT_B124 16'h9C3F
`define CUBE_LUT_B123 16'h9C3C
`define CUBE_LUT_B122 16'h9C3A
`define CUBE_LUT_B121 16'h9C37
`define CUBE_LUT_B120 16'h9C35
`define CUBE_LUT_B11F 16'h9C32
`define CUBE_LUT_B11E 16'h9C30
`define CUBE_LUT_B11D 16'h9C2E
`define CUBE_LUT_B11C 16'h9C2B
`define CUBE_LUT_B11B 16'h9C29
`define CUBE_LUT_B11A 16'h9C26
`define CUBE_LUT_B119 16'h9C24
`define CUBE_LUT_B118 16'h9C21
`define CUBE_LUT_B117 16'h9C1F
`define CUBE_LUT_B116 16'h9C1C
`define CUBE_LUT_B115 16'h9C1A
`define CUBE_LUT_B114 16'h9C18
`define CUBE_LUT_B113 16'h9C15
`define CUBE_LUT_B112 16'h9C13
`define CUBE_LUT_B111 16'h9C10
`define CUBE_LUT_B110 16'h9C0E
`define CUBE_LUT_B10F 16'h9C0C
`define CUBE_LUT_B10E 16'h9C09
`define CUBE_LUT_B10D 16'h9C07
`define CUBE_LUT_B10C 16'h9C04
`define CUBE_LUT_B10B 16'h9C02
`define CUBE_LUT_B10A 16'h9BFF
`define CUBE_LUT_B109 16'h9BFA
`define CUBE_LUT_B108 16'h9BF6
`define CUBE_LUT_B107 16'h9BF1
`define CUBE_LUT_B106 16'h9BEC
`define CUBE_LUT_B105 16'h9BE8
`define CUBE_LUT_B104 16'h9BE3
`define CUBE_LUT_B103 16'h9BDE
`define CUBE_LUT_B102 16'h9BD9
`define CUBE_LUT_B101 16'h9BD5
`define CUBE_LUT_B100 16'h9BD0
`define CUBE_LUT_B0FF 16'h9BCB
`define CUBE_LUT_B0FE 16'h9BC7
`define CUBE_LUT_B0FD 16'h9BC2
`define CUBE_LUT_B0FC 16'h9BBD
`define CUBE_LUT_B0FB 16'h9BB9
`define CUBE_LUT_B0FA 16'h9BB4
`define CUBE_LUT_B0F9 16'h9BAF
`define CUBE_LUT_B0F8 16'h9BAB
`define CUBE_LUT_B0F7 16'h9BA6
`define CUBE_LUT_B0F6 16'h9BA1
`define CUBE_LUT_B0F5 16'h9B9D
`define CUBE_LUT_B0F4 16'h9B98
`define CUBE_LUT_B0F3 16'h9B94
`define CUBE_LUT_B0F2 16'h9B8F
`define CUBE_LUT_B0F1 16'h9B8B
`define CUBE_LUT_B0F0 16'h9B86
`define CUBE_LUT_B0EF 16'h9B81
`define CUBE_LUT_B0EE 16'h9B7D
`define CUBE_LUT_B0ED 16'h9B78
`define CUBE_LUT_B0EC 16'h9B74
`define CUBE_LUT_B0EB 16'h9B6F
`define CUBE_LUT_B0EA 16'h9B6B
`define CUBE_LUT_B0E9 16'h9B66
`define CUBE_LUT_B0E8 16'h9B62
`define CUBE_LUT_B0E7 16'h9B5D
`define CUBE_LUT_B0E6 16'h9B59
`define CUBE_LUT_B0E5 16'h9B54
`define CUBE_LUT_B0E4 16'h9B50
`define CUBE_LUT_B0E3 16'h9B4B
`define CUBE_LUT_B0E2 16'h9B47
`define CUBE_LUT_B0E1 16'h9B42
`define CUBE_LUT_B0E0 16'h9B3E
`define CUBE_LUT_B0DF 16'h9B39
`define CUBE_LUT_B0DE 16'h9B35
`define CUBE_LUT_B0DD 16'h9B30
`define CUBE_LUT_B0DC 16'h9B2C
`define CUBE_LUT_B0DB 16'h9B28
`define CUBE_LUT_B0DA 16'h9B23
`define CUBE_LUT_B0D9 16'h9B1F
`define CUBE_LUT_B0D8 16'h9B1A
`define CUBE_LUT_B0D7 16'h9B16
`define CUBE_LUT_B0D6 16'h9B12
`define CUBE_LUT_B0D5 16'h9B0D
`define CUBE_LUT_B0D4 16'h9B09
`define CUBE_LUT_B0D3 16'h9B04
`define CUBE_LUT_B0D2 16'h9B00
`define CUBE_LUT_B0D1 16'h9AFC
`define CUBE_LUT_B0D0 16'h9AF7
`define CUBE_LUT_B0CF 16'h9AF3
`define CUBE_LUT_B0CE 16'h9AEF
`define CUBE_LUT_B0CD 16'h9AEA
`define CUBE_LUT_B0CC 16'h9AE6
`define CUBE_LUT_B0CB 16'h9AE2
`define CUBE_LUT_B0CA 16'h9ADD
`define CUBE_LUT_B0C9 16'h9AD9
`define CUBE_LUT_B0C8 16'h9AD5
`define CUBE_LUT_B0C7 16'h9AD1
`define CUBE_LUT_B0C6 16'h9ACC
`define CUBE_LUT_B0C5 16'h9AC8
`define CUBE_LUT_B0C4 16'h9AC4
`define CUBE_LUT_B0C3 16'h9ABF
`define CUBE_LUT_B0C2 16'h9ABB
`define CUBE_LUT_B0C1 16'h9AB7
`define CUBE_LUT_B0C0 16'h9AB3
`define CUBE_LUT_B0BF 16'h9AAF
`define CUBE_LUT_B0BE 16'h9AAA
`define CUBE_LUT_B0BD 16'h9AA6
`define CUBE_LUT_B0BC 16'h9AA2
`define CUBE_LUT_B0BB 16'h9A9E
`define CUBE_LUT_B0BA 16'h9A99
`define CUBE_LUT_B0B9 16'h9A95
`define CUBE_LUT_B0B8 16'h9A91
`define CUBE_LUT_B0B7 16'h9A8D
`define CUBE_LUT_B0B6 16'h9A89
`define CUBE_LUT_B0B5 16'h9A85
`define CUBE_LUT_B0B4 16'h9A80
`define CUBE_LUT_B0B3 16'h9A7C
`define CUBE_LUT_B0B2 16'h9A78
`define CUBE_LUT_B0B1 16'h9A74
`define CUBE_LUT_B0B0 16'h9A70
`define CUBE_LUT_B0AF 16'h9A6C
`define CUBE_LUT_B0AE 16'h9A68
`define CUBE_LUT_B0AD 16'h9A64
`define CUBE_LUT_B0AC 16'h9A60
`define CUBE_LUT_B0AB 16'h9A5B
`define CUBE_LUT_B0AA 16'h9A57
`define CUBE_LUT_B0A9 16'h9A53
`define CUBE_LUT_B0A8 16'h9A4F
`define CUBE_LUT_B0A7 16'h9A4B
`define CUBE_LUT_B0A6 16'h9A47
`define CUBE_LUT_B0A5 16'h9A43
`define CUBE_LUT_B0A4 16'h9A3F
`define CUBE_LUT_B0A3 16'h9A3B
`define CUBE_LUT_B0A2 16'h9A37
`define CUBE_LUT_B0A1 16'h9A33
`define CUBE_LUT_B0A0 16'h9A2F
`define CUBE_LUT_B09F 16'h9A2B
`define CUBE_LUT_B09E 16'h9A27
`define CUBE_LUT_B09D 16'h9A23
`define CUBE_LUT_B09C 16'h9A1F
`define CUBE_LUT_B09B 16'h9A1B
`define CUBE_LUT_B09A 16'h9A17
`define CUBE_LUT_B099 16'h9A13
`define CUBE_LUT_B098 16'h9A0F
`define CUBE_LUT_B097 16'h9A0B
`define CUBE_LUT_B096 16'h9A07
`define CUBE_LUT_B095 16'h9A03
`define CUBE_LUT_B094 16'h99FF
`define CUBE_LUT_B093 16'h99FB
`define CUBE_LUT_B092 16'h99F7
`define CUBE_LUT_B091 16'h99F4
`define CUBE_LUT_B090 16'h99F0
`define CUBE_LUT_B08F 16'h99EC
`define CUBE_LUT_B08E 16'h99E8
`define CUBE_LUT_B08D 16'h99E4
`define CUBE_LUT_B08C 16'h99E0
`define CUBE_LUT_B08B 16'h99DC
`define CUBE_LUT_B08A 16'h99D8
`define CUBE_LUT_B089 16'h99D4
`define CUBE_LUT_B088 16'h99D1
`define CUBE_LUT_B087 16'h99CD
`define CUBE_LUT_B086 16'h99C9
`define CUBE_LUT_B085 16'h99C5
`define CUBE_LUT_B084 16'h99C1
`define CUBE_LUT_B083 16'h99BD
`define CUBE_LUT_B082 16'h99BA
`define CUBE_LUT_B081 16'h99B6
`define CUBE_LUT_B080 16'h99B2
`define CUBE_LUT_B07F 16'h99AE
`define CUBE_LUT_B07E 16'h99AA
`define CUBE_LUT_B07D 16'h99A7
`define CUBE_LUT_B07C 16'h99A3
`define CUBE_LUT_B07B 16'h999F
`define CUBE_LUT_B07A 16'h999B
`define CUBE_LUT_B079 16'h9998
`define CUBE_LUT_B078 16'h9994
`define CUBE_LUT_B077 16'h9990
`define CUBE_LUT_B076 16'h998C
`define CUBE_LUT_B075 16'h9989
`define CUBE_LUT_B074 16'h9985
`define CUBE_LUT_B073 16'h9981
`define CUBE_LUT_B072 16'h997D
`define CUBE_LUT_B071 16'h997A
`define CUBE_LUT_B070 16'h9976
`define CUBE_LUT_B06F 16'h9972
`define CUBE_LUT_B06E 16'h996F
`define CUBE_LUT_B06D 16'h996B
`define CUBE_LUT_B06C 16'h9967
`define CUBE_LUT_B06B 16'h9964
`define CUBE_LUT_B06A 16'h9960
`define CUBE_LUT_B069 16'h995C
`define CUBE_LUT_B068 16'h9959
`define CUBE_LUT_B067 16'h9955
`define CUBE_LUT_B066 16'h9951
`define CUBE_LUT_B065 16'h994E
`define CUBE_LUT_B064 16'h994A
`define CUBE_LUT_B063 16'h9947
`define CUBE_LUT_B062 16'h9943
`define CUBE_LUT_B061 16'h993F
`define CUBE_LUT_B060 16'h993C
`define CUBE_LUT_B05F 16'h9938
`define CUBE_LUT_B05E 16'h9935
`define CUBE_LUT_B05D 16'h9931
`define CUBE_LUT_B05C 16'h992E
`define CUBE_LUT_B05B 16'h992A
`define CUBE_LUT_B05A 16'h9926
`define CUBE_LUT_B059 16'h9923
`define CUBE_LUT_B058 16'h991F
`define CUBE_LUT_B057 16'h991C
`define CUBE_LUT_B056 16'h9918
`define CUBE_LUT_B055 16'h9915
`define CUBE_LUT_B054 16'h9911
`define CUBE_LUT_B053 16'h990E
`define CUBE_LUT_B052 16'h990A
`define CUBE_LUT_B051 16'h9907
`define CUBE_LUT_B050 16'h9903
`define CUBE_LUT_B04F 16'h9900
`define CUBE_LUT_B04E 16'h98FC
`define CUBE_LUT_B04D 16'h98F9
`define CUBE_LUT_B04C 16'h98F5
`define CUBE_LUT_B04B 16'h98F2
`define CUBE_LUT_B04A 16'h98EE
`define CUBE_LUT_B049 16'h98EB
`define CUBE_LUT_B048 16'h98E8
`define CUBE_LUT_B047 16'h98E4
`define CUBE_LUT_B046 16'h98E1
`define CUBE_LUT_B045 16'h98DD
`define CUBE_LUT_B044 16'h98DA
`define CUBE_LUT_B043 16'h98D6
`define CUBE_LUT_B042 16'h98D3
`define CUBE_LUT_B041 16'h98D0
`define CUBE_LUT_B040 16'h98CC
`define CUBE_LUT_B03F 16'h98C9
`define CUBE_LUT_B03E 16'h98C5
`define CUBE_LUT_B03D 16'h98C2
`define CUBE_LUT_B03C 16'h98BF
`define CUBE_LUT_B03B 16'h98BB
`define CUBE_LUT_B03A 16'h98B8
`define CUBE_LUT_B039 16'h98B5
`define CUBE_LUT_B038 16'h98B1
`define CUBE_LUT_B037 16'h98AE
`define CUBE_LUT_B036 16'h98AB
`define CUBE_LUT_B035 16'h98A7
`define CUBE_LUT_B034 16'h98A4
`define CUBE_LUT_B033 16'h98A1
`define CUBE_LUT_B032 16'h989D
`define CUBE_LUT_B031 16'h989A
`define CUBE_LUT_B030 16'h9897
`define CUBE_LUT_B02F 16'h9894
`define CUBE_LUT_B02E 16'h9890
`define CUBE_LUT_B02D 16'h988D
`define CUBE_LUT_B02C 16'h988A
`define CUBE_LUT_B02B 16'h9886
`define CUBE_LUT_B02A 16'h9883
`define CUBE_LUT_B029 16'h9880
`define CUBE_LUT_B028 16'h987D
`define CUBE_LUT_B027 16'h987A
`define CUBE_LUT_B026 16'h9876
`define CUBE_LUT_B025 16'h9873
`define CUBE_LUT_B024 16'h9870
`define CUBE_LUT_B023 16'h986D
`define CUBE_LUT_B022 16'h9869
`define CUBE_LUT_B021 16'h9866
`define CUBE_LUT_B020 16'h9863
`define CUBE_LUT_B01F 16'h9860
`define CUBE_LUT_B01E 16'h985D
`define CUBE_LUT_B01D 16'h9859
`define CUBE_LUT_B01C 16'h9856
`define CUBE_LUT_B01B 16'h9853
`define CUBE_LUT_B01A 16'h9850
`define CUBE_LUT_B019 16'h984D
`define CUBE_LUT_B018 16'h984A
`define CUBE_LUT_B017 16'h9847
`define CUBE_LUT_B016 16'h9843
`define CUBE_LUT_B015 16'h9840
`define CUBE_LUT_B014 16'h983D
`define CUBE_LUT_B013 16'h983A
`define CUBE_LUT_B012 16'h9837
`define CUBE_LUT_B011 16'h9834
`define CUBE_LUT_B010 16'h9831
`define CUBE_LUT_B00F 16'h982E
`define CUBE_LUT_B00E 16'h982B
`define CUBE_LUT_B00D 16'h9827
`define CUBE_LUT_B00C 16'h9824
`define CUBE_LUT_B00B 16'h9821
`define CUBE_LUT_B00A 16'h981E
`define CUBE_LUT_B009 16'h981B
`define CUBE_LUT_B008 16'h9818
`define CUBE_LUT_B007 16'h9815
`define CUBE_LUT_B006 16'h9812
`define CUBE_LUT_B005 16'h980F
`define CUBE_LUT_B004 16'h980C
`define CUBE_LUT_B003 16'h9809
`define CUBE_LUT_B002 16'h9806
`define CUBE_LUT_B001 16'h9803
`define CUBE_LUT_B000 16'h9800
`define CUBE_LUT_AFFF 16'h97FD
`define CUBE_LUT_AFFD 16'h97F7
`define CUBE_LUT_AFFC 16'h97F4
`define CUBE_LUT_AFFB 16'h97F1
`define CUBE_LUT_AFFA 16'h97EE
`define CUBE_LUT_AFF8 16'h97E8
`define CUBE_LUT_AFF7 16'h97E5
`define CUBE_LUT_AFF6 16'h97E2
`define CUBE_LUT_AFF5 16'h97DF
`define CUBE_LUT_AFF4 16'h97DC
`define CUBE_LUT_AFF2 16'h97D6
`define CUBE_LUT_AFF1 16'h97D3
`define CUBE_LUT_AFF0 16'h97D0
`define CUBE_LUT_AFEF 16'h97CD
`define CUBE_LUT_AFED 16'h97C8
`define CUBE_LUT_AFEC 16'h97C5
`define CUBE_LUT_AFEB 16'h97C2
`define CUBE_LUT_AFEA 16'h97BF
`define CUBE_LUT_AFE8 16'h97B9
`define CUBE_LUT_AFE7 16'h97B6
`define CUBE_LUT_AFE6 16'h97B3
`define CUBE_LUT_AFE5 16'h97B0
`define CUBE_LUT_AFE4 16'h97AD
`define CUBE_LUT_AFE2 16'h97A7
`define CUBE_LUT_AFE1 16'h97A4
`define CUBE_LUT_AFE0 16'h97A1
`define CUBE_LUT_AFDF 16'h979F
`define CUBE_LUT_AFDD 16'h9799
`define CUBE_LUT_AFDC 16'h9796
`define CUBE_LUT_AFDB 16'h9793
`define CUBE_LUT_AFDA 16'h9790
`define CUBE_LUT_AFD8 16'h978A
`define CUBE_LUT_AFD7 16'h9787
`define CUBE_LUT_AFD6 16'h9785
`define CUBE_LUT_AFD5 16'h9782
`define CUBE_LUT_AFD4 16'h977F
`define CUBE_LUT_AFD2 16'h9779
`define CUBE_LUT_AFD1 16'h9776
`define CUBE_LUT_AFD0 16'h9773
`define CUBE_LUT_AFCF 16'h9770
`define CUBE_LUT_AFCD 16'h976B
`define CUBE_LUT_AFCC 16'h9768
`define CUBE_LUT_AFCB 16'h9765
`define CUBE_LUT_AFCA 16'h9762
`define CUBE_LUT_AFC9 16'h975F
`define CUBE_LUT_AFC7 16'h975A
`define CUBE_LUT_AFC6 16'h9757
`define CUBE_LUT_AFC5 16'h9754
`define CUBE_LUT_AFC4 16'h9751
`define CUBE_LUT_AFC2 16'h974C
`define CUBE_LUT_AFC1 16'h9749
`define CUBE_LUT_AFC0 16'h9746
`define CUBE_LUT_AFBF 16'h9743
`define CUBE_LUT_AFBD 16'h973E
`define CUBE_LUT_AFBC 16'h973B
`define CUBE_LUT_AFBB 16'h9738
`define CUBE_LUT_AFBA 16'h9735
`define CUBE_LUT_AFB9 16'h9732
`define CUBE_LUT_AFB7 16'h972D
`define CUBE_LUT_AFB6 16'h972A
`define CUBE_LUT_AFB5 16'h9727
`define CUBE_LUT_AFB4 16'h9724
`define CUBE_LUT_AFB2 16'h971F
`define CUBE_LUT_AFB1 16'h971C
`define CUBE_LUT_AFB0 16'h9719
`define CUBE_LUT_AFAF 16'h9716
`define CUBE_LUT_AFAD 16'h9711
`define CUBE_LUT_AFAC 16'h970E
`define CUBE_LUT_AFAB 16'h970B
`define CUBE_LUT_AFAA 16'h9709
`define CUBE_LUT_AFA9 16'h9706
`define CUBE_LUT_AFA7 16'h9700
`define CUBE_LUT_AFA6 16'h96FE
`define CUBE_LUT_AFA5 16'h96FB
`define CUBE_LUT_AFA4 16'h96F8
`define CUBE_LUT_AFA2 16'h96F3
`define CUBE_LUT_AFA1 16'h96F0
`define CUBE_LUT_AFA0 16'h96ED
`define CUBE_LUT_AF9F 16'h96EB
`define CUBE_LUT_AF9E 16'h96E8
`define CUBE_LUT_AF9C 16'h96E2
`define CUBE_LUT_AF9B 16'h96E0
`define CUBE_LUT_AF9A 16'h96DD
`define CUBE_LUT_AF99 16'h96DA
`define CUBE_LUT_AF97 16'h96D5
`define CUBE_LUT_AF96 16'h96D2
`define CUBE_LUT_AF95 16'h96CF
`define CUBE_LUT_AF94 16'h96CD
`define CUBE_LUT_AF92 16'h96C7
`define CUBE_LUT_AF91 16'h96C5
`define CUBE_LUT_AF90 16'h96C2
`define CUBE_LUT_AF8F 16'h96BF
`define CUBE_LUT_AF8E 16'h96BD
`define CUBE_LUT_AF8C 16'h96B7
`define CUBE_LUT_AF8B 16'h96B5
`define CUBE_LUT_AF8A 16'h96B2
`define CUBE_LUT_AF89 16'h96AF
`define CUBE_LUT_AF87 16'h96AA
`define CUBE_LUT_AF86 16'h96A7
`define CUBE_LUT_AF85 16'h96A5
`define CUBE_LUT_AF84 16'h96A2
`define CUBE_LUT_AF82 16'h969D
`define CUBE_LUT_AF81 16'h969A
`define CUBE_LUT_AF80 16'h9698
`define CUBE_LUT_AF7F 16'h9695
`define CUBE_LUT_AF7E 16'h9692
`define CUBE_LUT_AF7C 16'h968D
`define CUBE_LUT_AF7B 16'h968A
`define CUBE_LUT_AF7A 16'h9688
`define CUBE_LUT_AF79 16'h9685
`define CUBE_LUT_AF77 16'h9680
`define CUBE_LUT_AF76 16'h967D
`define CUBE_LUT_AF75 16'h967B
`define CUBE_LUT_AF74 16'h9678
`define CUBE_LUT_AF73 16'h9675
`define CUBE_LUT_AF71 16'h9670
`define CUBE_LUT_AF70 16'h966E
`define CUBE_LUT_AF6F 16'h966B
`define CUBE_LUT_AF6E 16'h9668
`define CUBE_LUT_AF6C 16'h9663
`define CUBE_LUT_AF6B 16'h9661
`define CUBE_LUT_AF6A 16'h965E
`define CUBE_LUT_AF69 16'h965C
`define CUBE_LUT_AF67 16'h9656
`define CUBE_LUT_AF66 16'h9654
`define CUBE_LUT_AF65 16'h9651
`define CUBE_LUT_AF64 16'h964F
`define CUBE_LUT_AF63 16'h964C
`define CUBE_LUT_AF61 16'h9647
`define CUBE_LUT_AF60 16'h9645
`define CUBE_LUT_AF5F 16'h9642
`define CUBE_LUT_AF5E 16'h963F
`define CUBE_LUT_AF5C 16'h963A
`define CUBE_LUT_AF5B 16'h9638
`define CUBE_LUT_AF5A 16'h9635
`define CUBE_LUT_AF59 16'h9633
`define CUBE_LUT_AF57 16'h962E
`define CUBE_LUT_AF56 16'h962B
`define CUBE_LUT_AF55 16'h9629
`define CUBE_LUT_AF54 16'h9626
`define CUBE_LUT_AF53 16'h9624
`define CUBE_LUT_AF51 16'h961F
`define CUBE_LUT_AF50 16'h961C
`define CUBE_LUT_AF4F 16'h961A
`define CUBE_LUT_AF4E 16'h9617
`define CUBE_LUT_AF4C 16'h9612
`define CUBE_LUT_AF4B 16'h9610
`define CUBE_LUT_AF4A 16'h960D
`define CUBE_LUT_AF49 16'h960B
`define CUBE_LUT_AF47 16'h9606
`define CUBE_LUT_AF46 16'h9603
`define CUBE_LUT_AF45 16'h9601
`define CUBE_LUT_AF44 16'h95FE
`define CUBE_LUT_AF43 16'h95FC
`define CUBE_LUT_AF41 16'h95F7
`define CUBE_LUT_AF40 16'h95F4
`define CUBE_LUT_AF3F 16'h95F2
`define CUBE_LUT_AF3E 16'h95EF
`define CUBE_LUT_AF3C 16'h95EA
`define CUBE_LUT_AF3B 16'h95E8
`define CUBE_LUT_AF3A 16'h95E6
`define CUBE_LUT_AF39 16'h95E3
`define CUBE_LUT_AF38 16'h95E1
`define CUBE_LUT_AF36 16'h95DC
`define CUBE_LUT_AF35 16'h95D9
`define CUBE_LUT_AF34 16'h95D7
`define CUBE_LUT_AF33 16'h95D5
`define CUBE_LUT_AF31 16'h95D0
`define CUBE_LUT_AF30 16'h95CD
`define CUBE_LUT_AF2F 16'h95CB
`define CUBE_LUT_AF2E 16'h95C8
`define CUBE_LUT_AF2C 16'h95C4
`define CUBE_LUT_AF2B 16'h95C1
`define CUBE_LUT_AF2A 16'h95BF
`define CUBE_LUT_AF29 16'h95BC
`define CUBE_LUT_AF28 16'h95BA
`define CUBE_LUT_AF26 16'h95B5
`define CUBE_LUT_AF25 16'h95B3
`define CUBE_LUT_AF24 16'h95B0
`define CUBE_LUT_AF23 16'h95AE
`define CUBE_LUT_AF21 16'h95A9
`define CUBE_LUT_AF20 16'h95A7
`define CUBE_LUT_AF1F 16'h95A4
`define CUBE_LUT_AF1E 16'h95A2
`define CUBE_LUT_AF1C 16'h959D
`define CUBE_LUT_AF1B 16'h959B
`define CUBE_LUT_AF1A 16'h9599
`define CUBE_LUT_AF19 16'h9596
`define CUBE_LUT_AF18 16'h9594
`define CUBE_LUT_AF16 16'h958F
`define CUBE_LUT_AF15 16'h958D
`define CUBE_LUT_AF14 16'h958A
`define CUBE_LUT_AF13 16'h9588
`define CUBE_LUT_AF11 16'h9583
`define CUBE_LUT_AF10 16'h9581
`define CUBE_LUT_AF0F 16'h957F
`define CUBE_LUT_AF0E 16'h957C
`define CUBE_LUT_AF0D 16'h957A
`define CUBE_LUT_AF0B 16'h9575
`define CUBE_LUT_AF0A 16'h9573
`define CUBE_LUT_AF09 16'h9571
`define CUBE_LUT_AF08 16'h956E
`define CUBE_LUT_AF06 16'h956A
`define CUBE_LUT_AF05 16'h9568
`define CUBE_LUT_AF04 16'h9565
`define CUBE_LUT_AF03 16'h9563
`define CUBE_LUT_AF01 16'h955E
`define CUBE_LUT_AF00 16'h955C
`define CUBE_LUT_AEFF 16'h955A
`define CUBE_LUT_AEFE 16'h9557
`define CUBE_LUT_AEFD 16'h9555
`define CUBE_LUT_AEFB 16'h9551
`define CUBE_LUT_AEFA 16'h954E
`define CUBE_LUT_AEF9 16'h954C
`define CUBE_LUT_AEF8 16'h954A
`define CUBE_LUT_AEF6 16'h9545
`define CUBE_LUT_AEF5 16'h9543
`define CUBE_LUT_AEF4 16'h9541
`define CUBE_LUT_AEF3 16'h953E
`define CUBE_LUT_AEF1 16'h953A
`define CUBE_LUT_AEF0 16'h9538
`define CUBE_LUT_AEEF 16'h9535
`define CUBE_LUT_AEEE 16'h9533
`define CUBE_LUT_AEED 16'h9531
`define CUBE_LUT_AEEB 16'h952C
`define CUBE_LUT_AEEA 16'h952A
`define CUBE_LUT_AEE9 16'h9528
`define CUBE_LUT_AEE8 16'h9526
`define CUBE_LUT_AEE6 16'h9521
`define CUBE_LUT_AEE5 16'h951F
`define CUBE_LUT_AEE4 16'h951D
`define CUBE_LUT_AEE3 16'h951A
`define CUBE_LUT_AEE2 16'h9518
`define CUBE_LUT_AEE0 16'h9514
`define CUBE_LUT_AEDF 16'h9512
`define CUBE_LUT_AEDE 16'h950F
`define CUBE_LUT_AEDD 16'h950D
`define CUBE_LUT_AEDB 16'h9509
`define CUBE_LUT_AEDA 16'h9507
`define CUBE_LUT_AED9 16'h9504
`define CUBE_LUT_AED8 16'h9502
`define CUBE_LUT_AED6 16'h94FE
`define CUBE_LUT_AED5 16'h94FC
`define CUBE_LUT_AED4 16'h94F9
`define CUBE_LUT_AED3 16'h94F7
`define CUBE_LUT_AED2 16'h94F5
`define CUBE_LUT_AED0 16'h94F1
`define CUBE_LUT_AECF 16'h94EF
`define CUBE_LUT_AECE 16'h94EC
`define CUBE_LUT_AECD 16'h94EA
`define CUBE_LUT_AECB 16'h94E6
`define CUBE_LUT_AECA 16'h94E4
`define CUBE_LUT_AEC9 16'h94E2
`define CUBE_LUT_AEC8 16'h94DF
`define CUBE_LUT_AEC6 16'h94DB
`define CUBE_LUT_AEC5 16'h94D9
`define CUBE_LUT_AEC4 16'h94D7
`define CUBE_LUT_AEC3 16'h94D5
`define CUBE_LUT_AEC2 16'h94D2
`define CUBE_LUT_AEC0 16'h94CE
`define CUBE_LUT_AEBF 16'h94CC
`define CUBE_LUT_AEBE 16'h94CA
`define CUBE_LUT_AEBD 16'h94C8
`define CUBE_LUT_AEBB 16'h94C4
`define CUBE_LUT_AEBA 16'h94C1
`define CUBE_LUT_AEB9 16'h94BF
`define CUBE_LUT_AEB8 16'h94BD
`define CUBE_LUT_AEB6 16'h94B9
`define CUBE_LUT_AEB5 16'h94B7
`define CUBE_LUT_AEB4 16'h94B5
`define CUBE_LUT_AEB3 16'h94B3
`define CUBE_LUT_AEB2 16'h94B1
`define CUBE_LUT_AEB0 16'h94AC
`define CUBE_LUT_AEAF 16'h94AA
`define CUBE_LUT_AEAE 16'h94A8
`define CUBE_LUT_AEAD 16'h94A6
`define CUBE_LUT_AEAB 16'h94A2
`define CUBE_LUT_AEAA 16'h94A0
`define CUBE_LUT_AEA9 16'h949E
`define CUBE_LUT_AEA8 16'h949C
`define CUBE_LUT_AEA7 16'h949A
`define CUBE_LUT_AEA5 16'h9495
`define CUBE_LUT_AEA4 16'h9493
`define CUBE_LUT_AEA3 16'h9491
`define CUBE_LUT_AEA2 16'h948F
`define CUBE_LUT_AEA0 16'h948B
`define CUBE_LUT_AE9F 16'h9489
`define CUBE_LUT_AE9E 16'h9487
`define CUBE_LUT_AE9D 16'h9485
`define CUBE_LUT_AE9B 16'h9481
`define CUBE_LUT_AE9A 16'h947F
`define CUBE_LUT_AE99 16'h947D
`define CUBE_LUT_AE98 16'h947B
`define CUBE_LUT_AE97 16'h9479
`define CUBE_LUT_AE95 16'h9475
`define CUBE_LUT_AE94 16'h9473
`define CUBE_LUT_AE93 16'h9471
`define CUBE_LUT_AE92 16'h946F
`define CUBE_LUT_AE90 16'h946A
`define CUBE_LUT_AE8F 16'h9468
`define CUBE_LUT_AE8E 16'h9466
`define CUBE_LUT_AE8D 16'h9464
`define CUBE_LUT_AE8B 16'h9460
`define CUBE_LUT_AE8A 16'h945E
`define CUBE_LUT_AE89 16'h945C
`define CUBE_LUT_AE88 16'h945A
`define CUBE_LUT_AE87 16'h9458
`define CUBE_LUT_AE85 16'h9454
`define CUBE_LUT_AE84 16'h9452
`define CUBE_LUT_AE83 16'h9450
`define CUBE_LUT_AE82 16'h944E
`define CUBE_LUT_AE80 16'h944A
`define CUBE_LUT_AE7F 16'h9449
`define CUBE_LUT_AE7E 16'h9447
`define CUBE_LUT_AE7D 16'h9445
`define CUBE_LUT_AE7C 16'h9443
`define CUBE_LUT_AE7A 16'h943F
`define CUBE_LUT_AE79 16'h943D
`define CUBE_LUT_AE78 16'h943B
`define CUBE_LUT_AE77 16'h9439
`define CUBE_LUT_AE75 16'h9435
`define CUBE_LUT_AE74 16'h9433
`define CUBE_LUT_AE73 16'h9431
`define CUBE_LUT_AE72 16'h942F
`define CUBE_LUT_AE70 16'h942B
`define CUBE_LUT_AE6F 16'h9429
`define CUBE_LUT_AE6E 16'h9427
`define CUBE_LUT_AE6D 16'h9425
`define CUBE_LUT_AE6C 16'h9423
`define CUBE_LUT_AE6A 16'h9420
`define CUBE_LUT_AE69 16'h941E
`define CUBE_LUT_AE68 16'h941C
`define CUBE_LUT_AE67 16'h941A
`define CUBE_LUT_AE65 16'h9416
`define CUBE_LUT_AE64 16'h9414
`define CUBE_LUT_AE63 16'h9412
`define CUBE_LUT_AE62 16'h9410
`define CUBE_LUT_AE60 16'h940C
`define CUBE_LUT_AE5F 16'h940A
`define CUBE_LUT_AE5E 16'h9409
`define CUBE_LUT_AE5D 16'h9407
`define CUBE_LUT_AE5C 16'h9405
`define CUBE_LUT_AE5A 16'h9401
`define CUBE_LUT_AE59 16'h93FE
`define CUBE_LUT_AE58 16'h93FA
`define CUBE_LUT_AE57 16'h93F7
`define CUBE_LUT_AE55 16'h93EF
`define CUBE_LUT_AE54 16'h93EB
`define CUBE_LUT_AE53 16'h93E8
`define CUBE_LUT_AE52 16'h93E4
`define CUBE_LUT_AE51 16'h93E0
`define CUBE_LUT_AE4F 16'h93D9
`define CUBE_LUT_AE4E 16'h93D5
`define CUBE_LUT_AE4D 16'h93D1
`define CUBE_LUT_AE4C 16'h93CD
`define CUBE_LUT_AE4A 16'h93C6
`define CUBE_LUT_AE49 16'h93C2
`define CUBE_LUT_AE48 16'h93BF
`define CUBE_LUT_AE47 16'h93BB
`define CUBE_LUT_AE45 16'h93B3
`define CUBE_LUT_AE44 16'h93B0
`define CUBE_LUT_AE43 16'h93AC
`define CUBE_LUT_AE42 16'h93A8
`define CUBE_LUT_AE41 16'h93A5
`define CUBE_LUT_AE3F 16'h939D
`define CUBE_LUT_AE3E 16'h939A
`define CUBE_LUT_AE3D 16'h9396
`define CUBE_LUT_AE3C 16'h9393
`define CUBE_LUT_AE3A 16'h938B
`define CUBE_LUT_AE39 16'h9388
`define CUBE_LUT_AE38 16'h9384
`define CUBE_LUT_AE37 16'h9380
`define CUBE_LUT_AE35 16'h9379
`define CUBE_LUT_AE34 16'h9376
`define CUBE_LUT_AE33 16'h9372
`define CUBE_LUT_AE32 16'h936E
`define CUBE_LUT_AE31 16'h936B
`define CUBE_LUT_AE2F 16'h9364
`define CUBE_LUT_AE2E 16'h9360
`define CUBE_LUT_AE2D 16'h935C
`define CUBE_LUT_AE2C 16'h9359
`define CUBE_LUT_AE2A 16'h9352
`define CUBE_LUT_AE29 16'h934E
`define CUBE_LUT_AE28 16'h934B
`define CUBE_LUT_AE27 16'h9347
`define CUBE_LUT_AE25 16'h9340
`define CUBE_LUT_AE24 16'h933C
`define CUBE_LUT_AE23 16'h9339
`define CUBE_LUT_AE22 16'h9335
`define CUBE_LUT_AE21 16'h9332
`define CUBE_LUT_AE1F 16'h932B
`define CUBE_LUT_AE1E 16'h9327
`define CUBE_LUT_AE1D 16'h9324
`define CUBE_LUT_AE1C 16'h9320
`define CUBE_LUT_AE1A 16'h9319
`define CUBE_LUT_AE19 16'h9316
`define CUBE_LUT_AE18 16'h9312
`define CUBE_LUT_AE17 16'h930F
`define CUBE_LUT_AE16 16'h930B
`define CUBE_LUT_AE14 16'h9304
`define CUBE_LUT_AE13 16'h9301
`define CUBE_LUT_AE12 16'h92FD
`define CUBE_LUT_AE11 16'h92FA
`define CUBE_LUT_AE0F 16'h92F3
`define CUBE_LUT_AE0E 16'h92F0
`define CUBE_LUT_AE0D 16'h92EC
`define CUBE_LUT_AE0C 16'h92E9
`define CUBE_LUT_AE0A 16'h92E2
`define CUBE_LUT_AE09 16'h92DF
`define CUBE_LUT_AE08 16'h92DB
`define CUBE_LUT_AE07 16'h92D8
`define CUBE_LUT_AE06 16'h92D4
`define CUBE_LUT_AE04 16'h92CE
`define CUBE_LUT_AE03 16'h92CA
`define CUBE_LUT_AE02 16'h92C7
`define CUBE_LUT_AE01 16'h92C3
`define CUBE_LUT_ADFF 16'h92BD
`define CUBE_LUT_ADFE 16'h92B9
`define CUBE_LUT_ADFD 16'h92B6
`define CUBE_LUT_ADFC 16'h92B3
`define CUBE_LUT_ADFA 16'h92AC
`define CUBE_LUT_ADF9 16'h92A8
`define CUBE_LUT_ADF8 16'h92A5
`define CUBE_LUT_ADF7 16'h92A2
`define CUBE_LUT_ADF6 16'h929E
`define CUBE_LUT_ADF4 16'h9298
`define CUBE_LUT_ADF3 16'h9294
`define CUBE_LUT_ADF2 16'h9291
`define CUBE_LUT_ADF1 16'h928E
`define CUBE_LUT_ADEF 16'h9287
`define CUBE_LUT_ADEE 16'h9284
`define CUBE_LUT_ADED 16'h9281
`define CUBE_LUT_ADEC 16'h927D
`define CUBE_LUT_ADEB 16'h927A
`define CUBE_LUT_ADE9 16'h9274
`define CUBE_LUT_ADE8 16'h9270
`define CUBE_LUT_ADE7 16'h926D
`define CUBE_LUT_ADE6 16'h926A
`define CUBE_LUT_ADE4 16'h9263
`define CUBE_LUT_ADE3 16'h9260
`define CUBE_LUT_ADE2 16'h925D
`define CUBE_LUT_ADE1 16'h9259
`define CUBE_LUT_ADDF 16'h9253
`define CUBE_LUT_ADDE 16'h9250
`define CUBE_LUT_ADDD 16'h924D
`define CUBE_LUT_ADDC 16'h9249
`define CUBE_LUT_ADDB 16'h9246
`define CUBE_LUT_ADD9 16'h9240
`define CUBE_LUT_ADD8 16'h923C
`define CUBE_LUT_ADD7 16'h9239
`define CUBE_LUT_ADD6 16'h9236
`define CUBE_LUT_ADD4 16'h9230
`define CUBE_LUT_ADD3 16'h922D
`define CUBE_LUT_ADD2 16'h9229
`define CUBE_LUT_ADD1 16'h9226
`define CUBE_LUT_ADCF 16'h9220
`define CUBE_LUT_ADCE 16'h921D
`define CUBE_LUT_ADCD 16'h921A
`define CUBE_LUT_ADCC 16'h9216
`define CUBE_LUT_ADCB 16'h9213
`define CUBE_LUT_ADC9 16'h920D
`define CUBE_LUT_ADC8 16'h920A
`define CUBE_LUT_ADC7 16'h9207
`define CUBE_LUT_ADC6 16'h9204
`define CUBE_LUT_ADC4 16'h91FD
`define CUBE_LUT_ADC3 16'h91FA
`define CUBE_LUT_ADC2 16'h91F7
`define CUBE_LUT_ADC1 16'h91F4
`define CUBE_LUT_ADC0 16'h91F1
`define CUBE_LUT_ADBE 16'h91EB
`define CUBE_LUT_ADBD 16'h91E8
`define CUBE_LUT_ADBC 16'h91E5
`define CUBE_LUT_ADBB 16'h91E1
`define CUBE_LUT_ADB9 16'h91DB
`define CUBE_LUT_ADB8 16'h91D8
`define CUBE_LUT_ADB7 16'h91D5
`define CUBE_LUT_ADB6 16'h91D2
`define CUBE_LUT_ADB4 16'h91CC
`define CUBE_LUT_ADB3 16'h91C9
`define CUBE_LUT_ADB2 16'h91C6
`define CUBE_LUT_ADB1 16'h91C3
`define CUBE_LUT_ADB0 16'h91C0
`define CUBE_LUT_ADAE 16'h91BA
`define CUBE_LUT_ADAD 16'h91B7
`define CUBE_LUT_ADAC 16'h91B4
`define CUBE_LUT_ADAB 16'h91B1
`define CUBE_LUT_ADA9 16'h91AB
`define CUBE_LUT_ADA8 16'h91A8
`define CUBE_LUT_ADA7 16'h91A5
`define CUBE_LUT_ADA6 16'h91A2
`define CUBE_LUT_ADA4 16'h919C
`define CUBE_LUT_ADA3 16'h9199
`define CUBE_LUT_ADA2 16'h9196
`define CUBE_LUT_ADA1 16'h9193
`define CUBE_LUT_ADA0 16'h9190
`define CUBE_LUT_AD9E 16'h918A
`define CUBE_LUT_AD9D 16'h9187
`define CUBE_LUT_AD9C 16'h9184
`define CUBE_LUT_AD9B 16'h9181
`define CUBE_LUT_AD99 16'h917B
`define CUBE_LUT_AD98 16'h9178
`define CUBE_LUT_AD97 16'h9175
`define CUBE_LUT_AD96 16'h9172
`define CUBE_LUT_AD94 16'h916D
`define CUBE_LUT_AD93 16'h916A
`define CUBE_LUT_AD92 16'h9167
`define CUBE_LUT_AD91 16'h9164
`define CUBE_LUT_AD90 16'h9161
`define CUBE_LUT_AD8E 16'h915B
`define CUBE_LUT_AD8D 16'h9158
`define CUBE_LUT_AD8C 16'h9155
`define CUBE_LUT_AD8B 16'h9152
`define CUBE_LUT_AD89 16'h914D
`define CUBE_LUT_AD88 16'h914A
`define CUBE_LUT_AD87 16'h9147
`define CUBE_LUT_AD86 16'h9144
`define CUBE_LUT_AD85 16'h9141
`define CUBE_LUT_AD83 16'h913C
`define CUBE_LUT_AD82 16'h9139
`define CUBE_LUT_AD81 16'h9136
`define CUBE_LUT_AD80 16'h9133
`define CUBE_LUT_AD7E 16'h912D
`define CUBE_LUT_AD7D 16'h912B
`define CUBE_LUT_AD7C 16'h9128
`define CUBE_LUT_AD7B 16'h9125
`define CUBE_LUT_AD79 16'h911F
`define CUBE_LUT_AD78 16'h911C
`define CUBE_LUT_AD77 16'h911A
`define CUBE_LUT_AD76 16'h9117
`define CUBE_LUT_AD75 16'h9114
`define CUBE_LUT_AD73 16'h910E
`define CUBE_LUT_AD72 16'h910C
`define CUBE_LUT_AD71 16'h9109
`define CUBE_LUT_AD70 16'h9106
`define CUBE_LUT_AD6E 16'h9101
`define CUBE_LUT_AD6D 16'h90FE
`define CUBE_LUT_AD6C 16'h90FB
`define CUBE_LUT_AD6B 16'h90F8
`define CUBE_LUT_AD69 16'h90F3
`define CUBE_LUT_AD68 16'h90F0
`define CUBE_LUT_AD67 16'h90ED
`define CUBE_LUT_AD66 16'h90EB
`define CUBE_LUT_AD65 16'h90E8
`define CUBE_LUT_AD63 16'h90E2
`define CUBE_LUT_AD62 16'h90E0
`define CUBE_LUT_AD61 16'h90DD
`define CUBE_LUT_AD60 16'h90DA
`define CUBE_LUT_AD5E 16'h90D5
`define CUBE_LUT_AD5D 16'h90D2
`define CUBE_LUT_AD5C 16'h90CF
`define CUBE_LUT_AD5B 16'h90CD
`define CUBE_LUT_AD5A 16'h90CA
`define CUBE_LUT_AD58 16'h90C5
`define CUBE_LUT_AD57 16'h90C2
`define CUBE_LUT_AD56 16'h90BF
`define CUBE_LUT_AD55 16'h90BD
`define CUBE_LUT_AD53 16'h90B7
`define CUBE_LUT_AD52 16'h90B5
`define CUBE_LUT_AD51 16'h90B2
`define CUBE_LUT_AD50 16'h90AF
`define CUBE_LUT_AD4E 16'h90AA
`define CUBE_LUT_AD4D 16'h90A8
`define CUBE_LUT_AD4C 16'h90A5
`define CUBE_LUT_AD4B 16'h90A2
`define CUBE_LUT_AD4A 16'h90A0
`define CUBE_LUT_AD48 16'h909A
`define CUBE_LUT_AD47 16'h9098
`define CUBE_LUT_AD46 16'h9095
`define CUBE_LUT_AD45 16'h9093
`define CUBE_LUT_AD43 16'h908D
`define CUBE_LUT_AD42 16'h908B
`define CUBE_LUT_AD41 16'h9088
`define CUBE_LUT_AD40 16'h9086
`define CUBE_LUT_AD3E 16'h9080
`define CUBE_LUT_AD3D 16'h907E
`define CUBE_LUT_AD3C 16'h907B
`define CUBE_LUT_AD3B 16'h9079
`define CUBE_LUT_AD3A 16'h9076
`define CUBE_LUT_AD38 16'h9071
`define CUBE_LUT_AD37 16'h906F
`define CUBE_LUT_AD36 16'h906C
`define CUBE_LUT_AD35 16'h9069
`define CUBE_LUT_AD33 16'h9064
`define CUBE_LUT_AD32 16'h9062
`define CUBE_LUT_AD31 16'h905F
`define CUBE_LUT_AD30 16'h905D
`define CUBE_LUT_AD2F 16'h905A
`define CUBE_LUT_AD2D 16'h9055
`define CUBE_LUT_AD2C 16'h9053
`define CUBE_LUT_AD2B 16'h9050
`define CUBE_LUT_AD2A 16'h904E
`define CUBE_LUT_AD28 16'h9049
`define CUBE_LUT_AD27 16'h9046
`define CUBE_LUT_AD26 16'h9044
`define CUBE_LUT_AD25 16'h9041
`define CUBE_LUT_AD23 16'h903C
`define CUBE_LUT_AD22 16'h903A
`define CUBE_LUT_AD21 16'h9037
`define CUBE_LUT_AD20 16'h9035
`define CUBE_LUT_AD1F 16'h9032
`define CUBE_LUT_AD1D 16'h902E
`define CUBE_LUT_AD1C 16'h902B
`define CUBE_LUT_AD1B 16'h9029
`define CUBE_LUT_AD1A 16'h9026
`define CUBE_LUT_AD18 16'h9021
`define CUBE_LUT_AD17 16'h901F
`define CUBE_LUT_AD16 16'h901C
`define CUBE_LUT_AD15 16'h901A
`define CUBE_LUT_AD13 16'h9015
`define CUBE_LUT_AD12 16'h9013
`define CUBE_LUT_AD11 16'h9010
`define CUBE_LUT_AD10 16'h900E
`define CUBE_LUT_AD0F 16'h900C
`define CUBE_LUT_AD0D 16'h9007
`define CUBE_LUT_AD0C 16'h9004
`define CUBE_LUT_AD0B 16'h9002
`define CUBE_LUT_AD0A 16'h8FFF
`define CUBE_LUT_AD08 16'h8FF6
`define CUBE_LUT_AD07 16'h8FF1
`define CUBE_LUT_AD06 16'h8FEC
`define CUBE_LUT_AD05 16'h8FE8
`define CUBE_LUT_AD03 16'h8FDE
`define CUBE_LUT_AD02 16'h8FD9
`define CUBE_LUT_AD01 16'h8FD5
`define CUBE_LUT_AD00 16'h8FD0
`define CUBE_LUT_ACFF 16'h8FCB
`define CUBE_LUT_ACFD 16'h8FC2
`define CUBE_LUT_ACFC 16'h8FBD
`define CUBE_LUT_ACFB 16'h8FB9
`define CUBE_LUT_ACFA 16'h8FB4
`define CUBE_LUT_ACF8 16'h8FAB
`define CUBE_LUT_ACF7 16'h8FA6
`define CUBE_LUT_ACF6 16'h8FA1
`define CUBE_LUT_ACF5 16'h8F9D
`define CUBE_LUT_ACF4 16'h8F98
`define CUBE_LUT_ACF2 16'h8F8F
`define CUBE_LUT_ACF1 16'h8F8B
`define CUBE_LUT_ACF0 16'h8F86
`define CUBE_LUT_ACEF 16'h8F81
`define CUBE_LUT_ACED 16'h8F78
`define CUBE_LUT_ACEC 16'h8F74
`define CUBE_LUT_ACEB 16'h8F6F
`define CUBE_LUT_ACEA 16'h8F6B
`define CUBE_LUT_ACE8 16'h8F62
`define CUBE_LUT_ACE7 16'h8F5D
`define CUBE_LUT_ACE6 16'h8F59
`define CUBE_LUT_ACE5 16'h8F54
`define CUBE_LUT_ACE4 16'h8F50
`define CUBE_LUT_ACE2 16'h8F47
`define CUBE_LUT_ACE1 16'h8F42
`define CUBE_LUT_ACE0 16'h8F3E
`define CUBE_LUT_ACDF 16'h8F39
`define CUBE_LUT_ACDD 16'h8F30
`define CUBE_LUT_ACDC 16'h8F2C
`define CUBE_LUT_ACDB 16'h8F28
`define CUBE_LUT_ACDA 16'h8F23
`define CUBE_LUT_ACD8 16'h8F1A
`define CUBE_LUT_ACD7 16'h8F16
`define CUBE_LUT_ACD6 16'h8F12
`define CUBE_LUT_ACD5 16'h8F0D
`define CUBE_LUT_ACD4 16'h8F09
`define CUBE_LUT_ACD2 16'h8F00
`define CUBE_LUT_ACD1 16'h8EFC
`define CUBE_LUT_ACD0 16'h8EF7
`define CUBE_LUT_ACCF 16'h8EF3
`define CUBE_LUT_ACCD 16'h8EEA
`define CUBE_LUT_ACCC 16'h8EE6
`define CUBE_LUT_ACCB 16'h8EE2
`define CUBE_LUT_ACCA 16'h8EDD
`define CUBE_LUT_ACC9 16'h8ED9
`define CUBE_LUT_ACC7 16'h8ED1
`define CUBE_LUT_ACC6 16'h8ECC
`define CUBE_LUT_ACC5 16'h8EC8
`define CUBE_LUT_ACC4 16'h8EC4
`define CUBE_LUT_ACC2 16'h8EBB
`define CUBE_LUT_ACC1 16'h8EB7
`define CUBE_LUT_ACC0 16'h8EB3
`define CUBE_LUT_ACBF 16'h8EAF
`define CUBE_LUT_ACBD 16'h8EA6
`define CUBE_LUT_ACBC 16'h8EA2
`define CUBE_LUT_ACBB 16'h8E9E
`define CUBE_LUT_ACBA 16'h8E99
`define CUBE_LUT_ACB9 16'h8E95
`define CUBE_LUT_ACB7 16'h8E8D
`define CUBE_LUT_ACB6 16'h8E89
`define CUBE_LUT_ACB5 16'h8E85
`define CUBE_LUT_ACB4 16'h8E80
`define CUBE_LUT_ACB2 16'h8E78
`define CUBE_LUT_ACB1 16'h8E74
`define CUBE_LUT_ACB0 16'h8E70
`define CUBE_LUT_ACAF 16'h8E6C
`define CUBE_LUT_ACAD 16'h8E64
`define CUBE_LUT_ACAC 16'h8E60
`define CUBE_LUT_ACAB 16'h8E5B
`define CUBE_LUT_ACAA 16'h8E57
`define CUBE_LUT_ACA9 16'h8E53
`define CUBE_LUT_ACA7 16'h8E4B
`define CUBE_LUT_ACA6 16'h8E47
`define CUBE_LUT_ACA5 16'h8E43
`define CUBE_LUT_ACA4 16'h8E3F
`define CUBE_LUT_ACA2 16'h8E37
`define CUBE_LUT_ACA1 16'h8E33
`define CUBE_LUT_ACA0 16'h8E2F
`define CUBE_LUT_AC9F 16'h8E2B
`define CUBE_LUT_AC9E 16'h8E27
`define CUBE_LUT_AC9C 16'h8E1F
`define CUBE_LUT_AC9B 16'h8E1B
`define CUBE_LUT_AC9A 16'h8E17
`define CUBE_LUT_AC99 16'h8E13
`define CUBE_LUT_AC97 16'h8E0B
`define CUBE_LUT_AC96 16'h8E07
`define CUBE_LUT_AC95 16'h8E03
`define CUBE_LUT_AC94 16'h8DFF
`define CUBE_LUT_AC92 16'h8DF7
`define CUBE_LUT_AC91 16'h8DF4
`define CUBE_LUT_AC90 16'h8DF0
`define CUBE_LUT_AC8F 16'h8DEC
`define CUBE_LUT_AC8E 16'h8DE8
`define CUBE_LUT_AC8C 16'h8DE0
`define CUBE_LUT_AC8B 16'h8DDC
`define CUBE_LUT_AC8A 16'h8DD8
`define CUBE_LUT_AC89 16'h8DD4
`define CUBE_LUT_AC87 16'h8DCD
`define CUBE_LUT_AC86 16'h8DC9
`define CUBE_LUT_AC85 16'h8DC5
`define CUBE_LUT_AC84 16'h8DC1
`define CUBE_LUT_AC82 16'h8DBA
`define CUBE_LUT_AC81 16'h8DB6
`define CUBE_LUT_AC80 16'h8DB2
`define CUBE_LUT_AC7F 16'h8DAE
`define CUBE_LUT_AC7E 16'h8DAA
`define CUBE_LUT_AC7C 16'h8DA3
`define CUBE_LUT_AC7B 16'h8D9F
`define CUBE_LUT_AC7A 16'h8D9B
`define CUBE_LUT_AC79 16'h8D98
`define CUBE_LUT_AC77 16'h8D90
`define CUBE_LUT_AC76 16'h8D8C
`define CUBE_LUT_AC75 16'h8D89
`define CUBE_LUT_AC74 16'h8D85
`define CUBE_LUT_AC72 16'h8D7D
`define CUBE_LUT_AC71 16'h8D7A
`define CUBE_LUT_AC70 16'h8D76
`define CUBE_LUT_AC6F 16'h8D72
`define CUBE_LUT_AC6E 16'h8D6F
`define CUBE_LUT_AC6C 16'h8D67
`define CUBE_LUT_AC6B 16'h8D64
`define CUBE_LUT_AC6A 16'h8D60
`define CUBE_LUT_AC69 16'h8D5C
`define CUBE_LUT_AC67 16'h8D55
`define CUBE_LUT_AC66 16'h8D51
`define CUBE_LUT_AC65 16'h8D4E
`define CUBE_LUT_AC64 16'h8D4A
`define CUBE_LUT_AC63 16'h8D47
`define CUBE_LUT_AC61 16'h8D3F
`define CUBE_LUT_AC60 16'h8D3C
`define CUBE_LUT_AC5F 16'h8D38
`define CUBE_LUT_AC5E 16'h8D35
`define CUBE_LUT_AC5C 16'h8D2E
`define CUBE_LUT_AC5B 16'h8D2A
`define CUBE_LUT_AC5A 16'h8D26
`define CUBE_LUT_AC59 16'h8D23
`define CUBE_LUT_AC57 16'h8D1C
`define CUBE_LUT_AC56 16'h8D18
`define CUBE_LUT_AC55 16'h8D15
`define CUBE_LUT_AC54 16'h8D11
`define CUBE_LUT_AC53 16'h8D0E
`define CUBE_LUT_AC51 16'h8D07
`define CUBE_LUT_AC50 16'h8D03
`define CUBE_LUT_AC4F 16'h8D00
`define CUBE_LUT_AC4E 16'h8CFC
`define CUBE_LUT_AC4C 16'h8CF5
`define CUBE_LUT_AC4B 16'h8CF2
`define CUBE_LUT_AC4A 16'h8CEE
`define CUBE_LUT_AC49 16'h8CEB
`define CUBE_LUT_AC47 16'h8CE4
`define CUBE_LUT_AC46 16'h8CE1
`define CUBE_LUT_AC45 16'h8CDD
`define CUBE_LUT_AC44 16'h8CDA
`define CUBE_LUT_AC43 16'h8CD6
`define CUBE_LUT_AC41 16'h8CD0
`define CUBE_LUT_AC40 16'h8CCC
`define CUBE_LUT_AC3F 16'h8CC9
`define CUBE_LUT_AC3E 16'h8CC5
`define CUBE_LUT_AC3C 16'h8CBF
`define CUBE_LUT_AC3B 16'h8CBB
`define CUBE_LUT_AC3A 16'h8CB8
`define CUBE_LUT_AC39 16'h8CB5
`define CUBE_LUT_AC38 16'h8CB1
`define CUBE_LUT_AC36 16'h8CAB
`define CUBE_LUT_AC35 16'h8CA7
`define CUBE_LUT_AC34 16'h8CA4
`define CUBE_LUT_AC33 16'h8CA1
`define CUBE_LUT_AC31 16'h8C9A
`define CUBE_LUT_AC30 16'h8C97
`define CUBE_LUT_AC2F 16'h8C94
`define CUBE_LUT_AC2E 16'h8C90
`define CUBE_LUT_AC2C 16'h8C8A
`define CUBE_LUT_AC2B 16'h8C86
`define CUBE_LUT_AC2A 16'h8C83
`define CUBE_LUT_AC29 16'h8C80
`define CUBE_LUT_AC28 16'h8C7D
`define CUBE_LUT_AC26 16'h8C76
`define CUBE_LUT_AC25 16'h8C73
`define CUBE_LUT_AC24 16'h8C70
`define CUBE_LUT_AC23 16'h8C6D
`define CUBE_LUT_AC21 16'h8C66
`define CUBE_LUT_AC20 16'h8C63
`define CUBE_LUT_AC1F 16'h8C60
`define CUBE_LUT_AC1E 16'h8C5D
`define CUBE_LUT_AC1C 16'h8C56
`define CUBE_LUT_AC1B 16'h8C53
`define CUBE_LUT_AC1A 16'h8C50
`define CUBE_LUT_AC19 16'h8C4D
`define CUBE_LUT_AC18 16'h8C4A
`define CUBE_LUT_AC16 16'h8C43
`define CUBE_LUT_AC15 16'h8C40
`define CUBE_LUT_AC14 16'h8C3D
`define CUBE_LUT_AC13 16'h8C3A
`define CUBE_LUT_AC11 16'h8C34
`define CUBE_LUT_AC10 16'h8C31
`define CUBE_LUT_AC0F 16'h8C2E
`define CUBE_LUT_AC0E 16'h8C2B
`define CUBE_LUT_AC0D 16'h8C27
`define CUBE_LUT_AC0B 16'h8C21
`define CUBE_LUT_AC0A 16'h8C1E
`define CUBE_LUT_AC09 16'h8C1B
`define CUBE_LUT_AC08 16'h8C18
`define CUBE_LUT_AC06 16'h8C12
`define CUBE_LUT_AC05 16'h8C0F
`define CUBE_LUT_AC04 16'h8C0C
`define CUBE_LUT_AC03 16'h8C09
`define CUBE_LUT_AC01 16'h8C03
`define CUBE_LUT_AC00 16'h8C00
`define CUBE_LUT_ABFE 16'h8BFA
`define CUBE_LUT_ABFC 16'h8BF4
`define CUBE_LUT_ABF9 16'h8BEB
`define CUBE_LUT_ABF7 16'h8BE5
`define CUBE_LUT_ABF4 16'h8BDC
`define CUBE_LUT_ABF2 16'h8BD6
`define CUBE_LUT_ABEF 16'h8BCD
`define CUBE_LUT_ABED 16'h8BC8
`define CUBE_LUT_ABEA 16'h8BBF
`define CUBE_LUT_ABE8 16'h8BB9
`define CUBE_LUT_ABE5 16'h8BB0
`define CUBE_LUT_ABE3 16'h8BAA
`define CUBE_LUT_ABE0 16'h8BA1
`define CUBE_LUT_ABDE 16'h8B9C
`define CUBE_LUT_ABDC 16'h8B96
`define CUBE_LUT_ABD9 16'h8B8D
`define CUBE_LUT_ABD7 16'h8B87
`define CUBE_LUT_ABD4 16'h8B7F
`define CUBE_LUT_ABD2 16'h8B79
`define CUBE_LUT_ABCF 16'h8B70
`define CUBE_LUT_ABCD 16'h8B6B
`define CUBE_LUT_ABCA 16'h8B62
`define CUBE_LUT_ABC8 16'h8B5D
`define CUBE_LUT_ABC5 16'h8B54
`define CUBE_LUT_ABC3 16'h8B4E
`define CUBE_LUT_ABC1 16'h8B49
`define CUBE_LUT_ABBE 16'h8B40
`define CUBE_LUT_ABBC 16'h8B3B
`define CUBE_LUT_ABB9 16'h8B32
`define CUBE_LUT_ABB7 16'h8B2D
`define CUBE_LUT_ABB4 16'h8B24
`define CUBE_LUT_ABB2 16'h8B1F
`define CUBE_LUT_ABAF 16'h8B16
`define CUBE_LUT_ABAD 16'h8B11
`define CUBE_LUT_ABAA 16'h8B09
`define CUBE_LUT_ABA8 16'h8B03
`define CUBE_LUT_ABA6 16'h8AFE
`define CUBE_LUT_ABA3 16'h8AF5
`define CUBE_LUT_ABA1 16'h8AF0
`define CUBE_LUT_AB9E 16'h8AE8
`define CUBE_LUT_AB9C 16'h8AE2
`define CUBE_LUT_AB99 16'h8ADA
`define CUBE_LUT_AB97 16'h8AD5
`define CUBE_LUT_AB94 16'h8ACD
`define CUBE_LUT_AB92 16'h8AC7
`define CUBE_LUT_AB8F 16'h8ABF
`define CUBE_LUT_AB8D 16'h8ABA
`define CUBE_LUT_AB8A 16'h8AB2
`define CUBE_LUT_AB88 16'h8AAD
`define CUBE_LUT_AB86 16'h8AA7
`define CUBE_LUT_AB83 16'h8A9F
`define CUBE_LUT_AB81 16'h8A9A
`define CUBE_LUT_AB7E 16'h8A92
`define CUBE_LUT_AB7C 16'h8A8D
`define CUBE_LUT_AB79 16'h8A85
`define CUBE_LUT_AB77 16'h8A80
`define CUBE_LUT_AB74 16'h8A78
`define CUBE_LUT_AB72 16'h8A73
`define CUBE_LUT_AB6F 16'h8A6B
`define CUBE_LUT_AB6D 16'h8A66
`define CUBE_LUT_AB6B 16'h8A61
`define CUBE_LUT_AB68 16'h8A59
`define CUBE_LUT_AB66 16'h8A54
`define CUBE_LUT_AB63 16'h8A4C
`define CUBE_LUT_AB61 16'h8A47
`define CUBE_LUT_AB5E 16'h8A3F
`define CUBE_LUT_AB5C 16'h8A3A
`define CUBE_LUT_AB59 16'h8A33
`define CUBE_LUT_AB57 16'h8A2E
`define CUBE_LUT_AB54 16'h8A26
`define CUBE_LUT_AB52 16'h8A21
`define CUBE_LUT_AB4F 16'h8A1A
`define CUBE_LUT_AB4D 16'h8A15
`define CUBE_LUT_AB4B 16'h8A10
`define CUBE_LUT_AB48 16'h8A08
`define CUBE_LUT_AB46 16'h8A03
`define CUBE_LUT_AB43 16'h89FC
`define CUBE_LUT_AB41 16'h89F7
`define CUBE_LUT_AB3E 16'h89EF
`define CUBE_LUT_AB3C 16'h89EA
`define CUBE_LUT_AB39 16'h89E3
`define CUBE_LUT_AB37 16'h89DE
`define CUBE_LUT_AB34 16'h89D7
`define CUBE_LUT_AB32 16'h89D2
`define CUBE_LUT_AB30 16'h89CD
`define CUBE_LUT_AB2D 16'h89C6
`define CUBE_LUT_AB2B 16'h89C1
`define CUBE_LUT_AB28 16'h89BA
`define CUBE_LUT_AB26 16'h89B5
`define CUBE_LUT_AB23 16'h89AE
`define CUBE_LUT_AB21 16'h89A9
`define CUBE_LUT_AB1E 16'h89A2
`define CUBE_LUT_AB1C 16'h899D
`define CUBE_LUT_AB19 16'h8996
`define CUBE_LUT_AB17 16'h8992
`define CUBE_LUT_AB15 16'h898D
`define CUBE_LUT_AB12 16'h8986
`define CUBE_LUT_AB10 16'h8981
`define CUBE_LUT_AB0D 16'h897A
`define CUBE_LUT_AB0B 16'h8975
`define CUBE_LUT_AB08 16'h896E
`define CUBE_LUT_AB06 16'h896A
`define CUBE_LUT_AB03 16'h8963
`define CUBE_LUT_AB01 16'h895E
`define CUBE_LUT_AAFE 16'h8957
`define CUBE_LUT_AAFC 16'h8953
`define CUBE_LUT_AAF9 16'h894C
`define CUBE_LUT_AAF7 16'h8947
`define CUBE_LUT_AAF5 16'h8943
`define CUBE_LUT_AAF2 16'h893C
`define CUBE_LUT_AAF0 16'h8938
`define CUBE_LUT_AAED 16'h8931
`define CUBE_LUT_AAEB 16'h892C
`define CUBE_LUT_AAE8 16'h8926
`define CUBE_LUT_AAE6 16'h8921
`define CUBE_LUT_AAE3 16'h891A
`define CUBE_LUT_AAE1 16'h8916
`define CUBE_LUT_AADE 16'h890F
`define CUBE_LUT_AADC 16'h890B
`define CUBE_LUT_AADA 16'h8907
`define CUBE_LUT_AAD7 16'h8900
`define CUBE_LUT_AAD5 16'h88FC
`define CUBE_LUT_AAD2 16'h88F5
`define CUBE_LUT_AAD0 16'h88F1
`define CUBE_LUT_AACD 16'h88EA
`define CUBE_LUT_AACB 16'h88E6
`define CUBE_LUT_AAC8 16'h88DF
`define CUBE_LUT_AAC6 16'h88DB
`define CUBE_LUT_AAC3 16'h88D5
`define CUBE_LUT_AAC1 16'h88D0
`define CUBE_LUT_AABE 16'h88CA
`define CUBE_LUT_AABC 16'h88C6
`define CUBE_LUT_AABA 16'h88C1
`define CUBE_LUT_AAB7 16'h88BB
`define CUBE_LUT_AAB5 16'h88B7
`define CUBE_LUT_AAB2 16'h88B1
`define CUBE_LUT_AAB0 16'h88AC
`define CUBE_LUT_AAAD 16'h88A6
`define CUBE_LUT_AAAB 16'h88A2
`define CUBE_LUT_AAA8 16'h889C
`define CUBE_LUT_AAA6 16'h8897
`define CUBE_LUT_AAA3 16'h8891
`define CUBE_LUT_AAA1 16'h888D
`define CUBE_LUT_AA9F 16'h8889
`define CUBE_LUT_AA9C 16'h8883
`define CUBE_LUT_AA9A 16'h887F
`define CUBE_LUT_AA97 16'h8879
`define CUBE_LUT_AA95 16'h8875
`define CUBE_LUT_AA92 16'h886F
`define CUBE_LUT_AA90 16'h886A
`define CUBE_LUT_AA8D 16'h8864
`define CUBE_LUT_AA8B 16'h8860
`define CUBE_LUT_AA88 16'h885A
`define CUBE_LUT_AA86 16'h8856
`define CUBE_LUT_AA84 16'h8852
`define CUBE_LUT_AA81 16'h884C
`define CUBE_LUT_AA7F 16'h8849
`define CUBE_LUT_AA7C 16'h8843
`define CUBE_LUT_AA7A 16'h883F
`define CUBE_LUT_AA77 16'h8839
`define CUBE_LUT_AA75 16'h8835
`define CUBE_LUT_AA72 16'h882F
`define CUBE_LUT_AA70 16'h882B
`define CUBE_LUT_AA6D 16'h8825
`define CUBE_LUT_AA6B 16'h8821
`define CUBE_LUT_AA68 16'h881C
`define CUBE_LUT_AA66 16'h8818
`define CUBE_LUT_AA64 16'h8814
`define CUBE_LUT_AA61 16'h880E
`define CUBE_LUT_AA5F 16'h880A
`define CUBE_LUT_AA5C 16'h8805
`define CUBE_LUT_AA5A 16'h8801
`define CUBE_LUT_AA57 16'h87F7
`define CUBE_LUT_AA55 16'h87EF
`define CUBE_LUT_AA52 16'h87E4
`define CUBE_LUT_AA50 16'h87DC
`define CUBE_LUT_AA4D 16'h87D1
`define CUBE_LUT_AA4B 16'h87CA
`define CUBE_LUT_AA49 16'h87C2
`define CUBE_LUT_AA46 16'h87B7
`define CUBE_LUT_AA44 16'h87B0
`define CUBE_LUT_AA41 16'h87A5
`define CUBE_LUT_AA3F 16'h879D
`define CUBE_LUT_AA3C 16'h8793
`define CUBE_LUT_AA3A 16'h878B
`define CUBE_LUT_AA37 16'h8780
`define CUBE_LUT_AA35 16'h8779
`define CUBE_LUT_AA32 16'h876E
`define CUBE_LUT_AA30 16'h8767
`define CUBE_LUT_AA2D 16'h875C
`define CUBE_LUT_AA2B 16'h8755
`define CUBE_LUT_AA29 16'h874E
`define CUBE_LUT_AA26 16'h8743
`define CUBE_LUT_AA24 16'h873C
`define CUBE_LUT_AA21 16'h8732
`define CUBE_LUT_AA1F 16'h872B
`define CUBE_LUT_AA1C 16'h8720
`define CUBE_LUT_AA1A 16'h8719
`define CUBE_LUT_AA17 16'h870F
`define CUBE_LUT_AA15 16'h8708
`define CUBE_LUT_AA12 16'h86FD
`define CUBE_LUT_AA10 16'h86F7
`define CUBE_LUT_AA0E 16'h86F0
`define CUBE_LUT_AA0B 16'h86E5
`define CUBE_LUT_AA09 16'h86DF
`define CUBE_LUT_AA06 16'h86D4
`define CUBE_LUT_AA04 16'h86CE
`define CUBE_LUT_AA01 16'h86C3
`define CUBE_LUT_A9FF 16'h86BD
`define CUBE_LUT_A9FC 16'h86B3
`define CUBE_LUT_A9FA 16'h86AC
`define CUBE_LUT_A9F7 16'h86A2
`define CUBE_LUT_A9F5 16'h869B
`define CUBE_LUT_A9F3 16'h8694
`define CUBE_LUT_A9F0 16'h868B
`define CUBE_LUT_A9EE 16'h8684
`define CUBE_LUT_A9EB 16'h867A
`define CUBE_LUT_A9E9 16'h8674
`define CUBE_LUT_A9E6 16'h866A
`define CUBE_LUT_A9E4 16'h8663
`define CUBE_LUT_A9E1 16'h8659
`define CUBE_LUT_A9DF 16'h8653
`define CUBE_LUT_A9DC 16'h8649
`define CUBE_LUT_A9DA 16'h8643
`define CUBE_LUT_A9D7 16'h8639
`define CUBE_LUT_A9D5 16'h8633
`define CUBE_LUT_A9D3 16'h862D
`define CUBE_LUT_A9D0 16'h8623
`define CUBE_LUT_A9CE 16'h861D
`define CUBE_LUT_A9CB 16'h8613
`define CUBE_LUT_A9C9 16'h860D
`define CUBE_LUT_A9C6 16'h8604
`define CUBE_LUT_A9C4 16'h85FD
`define CUBE_LUT_A9C1 16'h85F4
`define CUBE_LUT_A9BF 16'h85EE
`define CUBE_LUT_A9BC 16'h85E5
`define CUBE_LUT_A9BA 16'h85DE
`define CUBE_LUT_A9B8 16'h85D8
`define CUBE_LUT_A9B5 16'h85CF
`define CUBE_LUT_A9B3 16'h85C9
`define CUBE_LUT_A9B0 16'h85C0
`define CUBE_LUT_A9AE 16'h85BA
`define CUBE_LUT_A9AB 16'h85B1
`define CUBE_LUT_A9A9 16'h85AB
`define CUBE_LUT_A9A6 16'h85A2
`define CUBE_LUT_A9A4 16'h859C
`define CUBE_LUT_A9A1 16'h8593
`define CUBE_LUT_A99F 16'h858D
`define CUBE_LUT_A99C 16'h8584
`define CUBE_LUT_A99A 16'h857E
`define CUBE_LUT_A998 16'h8578
`define CUBE_LUT_A995 16'h856F
`define CUBE_LUT_A993 16'h856A
`define CUBE_LUT_A990 16'h8561
`define CUBE_LUT_A98E 16'h855B
`define CUBE_LUT_A98B 16'h8552
`define CUBE_LUT_A989 16'h854D
`define CUBE_LUT_A986 16'h8544
`define CUBE_LUT_A984 16'h853E
`define CUBE_LUT_A981 16'h8536
`define CUBE_LUT_A97F 16'h8530
`define CUBE_LUT_A97D 16'h852B
`define CUBE_LUT_A97A 16'h8522
`define CUBE_LUT_A978 16'h851C
`define CUBE_LUT_A975 16'h8514
`define CUBE_LUT_A973 16'h850E
`define CUBE_LUT_A970 16'h8506
`define CUBE_LUT_A96E 16'h8501
`define CUBE_LUT_A96B 16'h84F8
`define CUBE_LUT_A969 16'h84F3
`define CUBE_LUT_A966 16'h84EB
`define CUBE_LUT_A964 16'h84E5
`define CUBE_LUT_A962 16'h84E0
`define CUBE_LUT_A95F 16'h84D8
`define CUBE_LUT_A95D 16'h84D2
`define CUBE_LUT_A95A 16'h84CA
`define CUBE_LUT_A958 16'h84C5
`define CUBE_LUT_A955 16'h84BD
`define CUBE_LUT_A953 16'h84B7
`define CUBE_LUT_A950 16'h84AF
`define CUBE_LUT_A94E 16'h84AA
`define CUBE_LUT_A94B 16'h84A2
`define CUBE_LUT_A949 16'h849D
`define CUBE_LUT_A946 16'h8495
`define CUBE_LUT_A944 16'h8490
`define CUBE_LUT_A942 16'h848B
`define CUBE_LUT_A93F 16'h8483
`define CUBE_LUT_A93D 16'h847E
`define CUBE_LUT_A93A 16'h8476
`define CUBE_LUT_A938 16'h8471
`define CUBE_LUT_A935 16'h8469
`define CUBE_LUT_A933 16'h8464
`define CUBE_LUT_A930 16'h845D
`define CUBE_LUT_A92E 16'h8458
`define CUBE_LUT_A92B 16'h8450
`define CUBE_LUT_A929 16'h844B
`define CUBE_LUT_A927 16'h8446
`define CUBE_LUT_A924 16'h843F
`define CUBE_LUT_A922 16'h843A
`define CUBE_LUT_A91F 16'h8432
`define CUBE_LUT_A91D 16'h842E
`define CUBE_LUT_A91A 16'h8426
`define CUBE_LUT_A918 16'h8421
`define CUBE_LUT_A915 16'h841A
`define CUBE_LUT_A913 16'h8415
`define CUBE_LUT_A910 16'h840E
`define CUBE_LUT_A90E 16'h8409
`define CUBE_LUT_A90B 16'h8402
`define CUBE_LUT_A909 16'h83FD
`define CUBE_LUT_A907 16'h83F8
`define CUBE_LUT_A904 16'h83F1
`define CUBE_LUT_A902 16'h83ED
`define CUBE_LUT_A8FF 16'h83E6
`define CUBE_LUT_A8FD 16'h83E1
`define CUBE_LUT_A8FA 16'h83DA
`define CUBE_LUT_A8F8 16'h83D5
`define CUBE_LUT_A8F5 16'h83CE
`define CUBE_LUT_A8F3 16'h83CA
`define CUBE_LUT_A8F0 16'h83C3
`define CUBE_LUT_A8EE 16'h83BE
`define CUBE_LUT_A8EC 16'h83BA
`define CUBE_LUT_A8E9 16'h83B3
`define CUBE_LUT_A8E7 16'h83AF
`define CUBE_LUT_A8E4 16'h83A8
`define CUBE_LUT_A8E2 16'h83A3
`define CUBE_LUT_A8DF 16'h839D
`define CUBE_LUT_A8DD 16'h8398
`define CUBE_LUT_A8DA 16'h8392
`define CUBE_LUT_A8D8 16'h838D
`define CUBE_LUT_A8D5 16'h8387
`define CUBE_LUT_A8D3 16'h8382
`define CUBE_LUT_A8D1 16'h837E
`define CUBE_LUT_A8CE 16'h8377
`define CUBE_LUT_A8CC 16'h8373
`define CUBE_LUT_A8C9 16'h836D
`define CUBE_LUT_A8C7 16'h8368
`define CUBE_LUT_A8C4 16'h8362
`define CUBE_LUT_A8C2 16'h835E
`define CUBE_LUT_A8BF 16'h8357
`define CUBE_LUT_A8BD 16'h8353
`define CUBE_LUT_A8BA 16'h834D
`define CUBE_LUT_A8B8 16'h8349
`define CUBE_LUT_A8B5 16'h8342
`define CUBE_LUT_A8B3 16'h833E
`define CUBE_LUT_A8B1 16'h833A
`define CUBE_LUT_A8AE 16'h8334
`define CUBE_LUT_A8AC 16'h8330
`define CUBE_LUT_A8A9 16'h832A
`define CUBE_LUT_A8A7 16'h8326
`define CUBE_LUT_A8A4 16'h8320
`define CUBE_LUT_A8A2 16'h831B
`define CUBE_LUT_A89F 16'h8315
`define CUBE_LUT_A89D 16'h8311
`define CUBE_LUT_A89A 16'h830B
`define CUBE_LUT_A898 16'h8308
`define CUBE_LUT_A896 16'h8304
`define CUBE_LUT_A893 16'h82FE
`define CUBE_LUT_A891 16'h82FA
`define CUBE_LUT_A88E 16'h82F4
`define CUBE_LUT_A88C 16'h82F0
`define CUBE_LUT_A889 16'h82EA
`define CUBE_LUT_A887 16'h82E6
`define CUBE_LUT_A884 16'h82E1
`define CUBE_LUT_A882 16'h82DD
`define CUBE_LUT_A87F 16'h82D7
`define CUBE_LUT_A87D 16'h82D3
`define CUBE_LUT_A87A 16'h82CE
`define CUBE_LUT_A878 16'h82CA
`define CUBE_LUT_A876 16'h82C6
`define CUBE_LUT_A873 16'h82C1
`define CUBE_LUT_A871 16'h82BD
`define CUBE_LUT_A86E 16'h82B7
`define CUBE_LUT_A86C 16'h82B4
`define CUBE_LUT_A869 16'h82AE
`define CUBE_LUT_A867 16'h82AB
`define CUBE_LUT_A864 16'h82A5
`define CUBE_LUT_A862 16'h82A2
`define CUBE_LUT_A85F 16'h829C
`define CUBE_LUT_A85D 16'h8299
`define CUBE_LUT_A85B 16'h8295
`define CUBE_LUT_A858 16'h8290
`define CUBE_LUT_A856 16'h828C
`define CUBE_LUT_A853 16'h8287
`define CUBE_LUT_A851 16'h8283
`define CUBE_LUT_A84E 16'h827E
`define CUBE_LUT_A84C 16'h827B
`define CUBE_LUT_A849 16'h8275
`define CUBE_LUT_A847 16'h8272
`define CUBE_LUT_A844 16'h826D
`define CUBE_LUT_A842 16'h826A
`define CUBE_LUT_A840 16'h8266
`define CUBE_LUT_A83D 16'h8261
`define CUBE_LUT_A83B 16'h825E
`define CUBE_LUT_A838 16'h8259
`define CUBE_LUT_A836 16'h8255
`define CUBE_LUT_A833 16'h8250
`define CUBE_LUT_A831 16'h824D
`define CUBE_LUT_A82E 16'h8248
`define CUBE_LUT_A82C 16'h8245
`define CUBE_LUT_A829 16'h8240
`define CUBE_LUT_A827 16'h823D
`define CUBE_LUT_A824 16'h8238
`define CUBE_LUT_A822 16'h8235
`define CUBE_LUT_A820 16'h8232
`define CUBE_LUT_A81D 16'h822D
`define CUBE_LUT_A81B 16'h822A
`define CUBE_LUT_A818 16'h8225
`define CUBE_LUT_A816 16'h8222
`define CUBE_LUT_A813 16'h821D
`define CUBE_LUT_A811 16'h821A
`define CUBE_LUT_A80E 16'h8215
`define CUBE_LUT_A80C 16'h8212
`define CUBE_LUT_A809 16'h820E
`define CUBE_LUT_A807 16'h820B
`define CUBE_LUT_A805 16'h8208
`define CUBE_LUT_A802 16'h8203
`define CUBE_LUT_A7FF 16'h81FF
`define CUBE_LUT_A7FA 16'h81FC
`define CUBE_LUT_A7F5 16'h81F8
`define CUBE_LUT_A7F0 16'h81F4
`define CUBE_LUT_A7EC 16'h81F1
`define CUBE_LUT_A7E7 16'h81ED
`define CUBE_LUT_A7E2 16'h81EA
`define CUBE_LUT_A7DD 16'h81E6
`define CUBE_LUT_A7D8 16'h81E3
`define CUBE_LUT_A7D3 16'h81DF
`define CUBE_LUT_A7CE 16'h81DB
`define CUBE_LUT_A7C9 16'h81D8
`define CUBE_LUT_A7C4 16'h81D4
`define CUBE_LUT_A7BF 16'h81D1
`define CUBE_LUT_A7BA 16'h81CD
`define CUBE_LUT_A7B5 16'h81CA
`define CUBE_LUT_A7B1 16'h81C7
`define CUBE_LUT_A7AC 16'h81C4
`define CUBE_LUT_A7A7 16'h81C0
`define CUBE_LUT_A7A2 16'h81BD
`define CUBE_LUT_A79D 16'h81B9
`define CUBE_LUT_A798 16'h81B6
`define CUBE_LUT_A793 16'h81B3
`define CUBE_LUT_A78E 16'h81AF
`define CUBE_LUT_A789 16'h81AC
`define CUBE_LUT_A784 16'h81A9
`define CUBE_LUT_A77F 16'h81A5
`define CUBE_LUT_A77A 16'h81A2
`define CUBE_LUT_A776 16'h819F
`define CUBE_LUT_A771 16'h819C
`define CUBE_LUT_A76C 16'h8199
`define CUBE_LUT_A767 16'h8196
`define CUBE_LUT_A762 16'h8192
`define CUBE_LUT_A75D 16'h818F
`define CUBE_LUT_A758 16'h818C
`define CUBE_LUT_A753 16'h8189
`define CUBE_LUT_A74E 16'h8186
`define CUBE_LUT_A749 16'h8183
`define CUBE_LUT_A744 16'h8180
`define CUBE_LUT_A740 16'h817D
`define CUBE_LUT_A73B 16'h817A
`define CUBE_LUT_A736 16'h8177
`define CUBE_LUT_A731 16'h8174
`define CUBE_LUT_A72C 16'h8171
`define CUBE_LUT_A727 16'h816E
`define CUBE_LUT_A722 16'h816B
`define CUBE_LUT_A71D 16'h8168
`define CUBE_LUT_A718 16'h8165
`define CUBE_LUT_A713 16'h8162
`define CUBE_LUT_A70E 16'h815F
`define CUBE_LUT_A709 16'h815C
`define CUBE_LUT_A705 16'h815A
`define CUBE_LUT_A700 16'h8157
`define CUBE_LUT_A6FB 16'h8154
`define CUBE_LUT_A6F6 16'h8151
`define CUBE_LUT_A6F1 16'h814E
`define CUBE_LUT_A6EC 16'h814C
`define CUBE_LUT_A6E7 16'h8149
`define CUBE_LUT_A6E2 16'h8146
`define CUBE_LUT_A6DD 16'h8143
`define CUBE_LUT_A6D8 16'h8141
`define CUBE_LUT_A6D3 16'h813E
`define CUBE_LUT_A6CE 16'h813B
`define CUBE_LUT_A6CA 16'h8139
`define CUBE_LUT_A6C5 16'h8136
`define CUBE_LUT_A6C0 16'h8134
`define CUBE_LUT_A6BB 16'h8131
`define CUBE_LUT_A6B6 16'h812E
`define CUBE_LUT_A6B1 16'h812C
`define CUBE_LUT_A6AC 16'h8129
`define CUBE_LUT_A6A7 16'h8126
`define CUBE_LUT_A6A2 16'h8124
`define CUBE_LUT_A69D 16'h8121
`define CUBE_LUT_A698 16'h811F
`define CUBE_LUT_A693 16'h811C
`define CUBE_LUT_A68F 16'h811A
`define CUBE_LUT_A68A 16'h8118
`define CUBE_LUT_A685 16'h8115
`define CUBE_LUT_A680 16'h8113
`define CUBE_LUT_A67B 16'h8110
`define CUBE_LUT_A676 16'h810E
`define CUBE_LUT_A671 16'h810B
`define CUBE_LUT_A66C 16'h8109
`define CUBE_LUT_A667 16'h8106
`define CUBE_LUT_A662 16'h8104
`define CUBE_LUT_A65D 16'h8102
`define CUBE_LUT_A658 16'h80FF
`define CUBE_LUT_A654 16'h80FD
`define CUBE_LUT_A64F 16'h80FB
`define CUBE_LUT_A64A 16'h80F9
`define CUBE_LUT_A645 16'h80F6
`define CUBE_LUT_A640 16'h80F4
`define CUBE_LUT_A63B 16'h80F2
`define CUBE_LUT_A636 16'h80F0
`define CUBE_LUT_A631 16'h80ED
`define CUBE_LUT_A62C 16'h80EB
`define CUBE_LUT_A627 16'h80E9
`define CUBE_LUT_A622 16'h80E7
`define CUBE_LUT_A61E 16'h80E5
`define CUBE_LUT_A619 16'h80E3
`define CUBE_LUT_A614 16'h80E1
`define CUBE_LUT_A60F 16'h80DE
`define CUBE_LUT_A60A 16'h80DC
`define CUBE_LUT_A605 16'h80DA
`define CUBE_LUT_A600 16'h80D8
`define CUBE_LUT_A5FB 16'h80D6
`define CUBE_LUT_A5F6 16'h80D4
`define CUBE_LUT_A5F1 16'h80D2
`define CUBE_LUT_A5EC 16'h80D0
`define CUBE_LUT_A5E7 16'h80CE
`define CUBE_LUT_A5E3 16'h80CC
`define CUBE_LUT_A5DE 16'h80CA
`define CUBE_LUT_A5D9 16'h80C8
`define CUBE_LUT_A5D4 16'h80C6
`define CUBE_LUT_A5CF 16'h80C4
`define CUBE_LUT_A5CA 16'h80C2
`define CUBE_LUT_A5C5 16'h80C0
`define CUBE_LUT_A5C0 16'h80BE
`define CUBE_LUT_A5BB 16'h80BC
`define CUBE_LUT_A5B6 16'h80BA
`define CUBE_LUT_A5B1 16'h80B8
`define CUBE_LUT_A5AC 16'h80B6
`define CUBE_LUT_A5A8 16'h80B5
`define CUBE_LUT_A5A3 16'h80B3
`define CUBE_LUT_A59E 16'h80B1
`define CUBE_LUT_A599 16'h80AF
`define CUBE_LUT_A594 16'h80AE
`define CUBE_LUT_A58F 16'h80AC
`define CUBE_LUT_A58A 16'h80AA
`define CUBE_LUT_A585 16'h80A8
`define CUBE_LUT_A580 16'h80A6
`define CUBE_LUT_A57B 16'h80A5
`define CUBE_LUT_A576 16'h80A3
`define CUBE_LUT_A571 16'h80A1
`define CUBE_LUT_A56D 16'h80A0
`define CUBE_LUT_A568 16'h809E
`define CUBE_LUT_A563 16'h809C
`define CUBE_LUT_A55E 16'h809B
`define CUBE_LUT_A559 16'h8099
`define CUBE_LUT_A554 16'h8097
`define CUBE_LUT_A54F 16'h8096
`define CUBE_LUT_A54A 16'h8094
`define CUBE_LUT_A545 16'h8092
`define CUBE_LUT_A540 16'h8091
`define CUBE_LUT_A53B 16'h808F
`define CUBE_LUT_A536 16'h808D
`define CUBE_LUT_A532 16'h808C
`define CUBE_LUT_A52D 16'h808B
`define CUBE_LUT_A528 16'h8089
`define CUBE_LUT_A523 16'h8088
`define CUBE_LUT_A51E 16'h8086
`define CUBE_LUT_A519 16'h8084
`define CUBE_LUT_A514 16'h8083
`define CUBE_LUT_A50F 16'h8081
`define CUBE_LUT_A50A 16'h8080
`define CUBE_LUT_A505 16'h807E
`define CUBE_LUT_A500 16'h807D
`define CUBE_LUT_A4FC 16'h807C
`define CUBE_LUT_A4F7 16'h807A
`define CUBE_LUT_A4F2 16'h8079
`define CUBE_LUT_A4ED 16'h8078
`define CUBE_LUT_A4E8 16'h8076
`define CUBE_LUT_A4E3 16'h8075
`define CUBE_LUT_A4DE 16'h8073
`define CUBE_LUT_A4D9 16'h8072
`define CUBE_LUT_A4D4 16'h8071
`define CUBE_LUT_A4CF 16'h806F
`define CUBE_LUT_A4CA 16'h806E
`define CUBE_LUT_A4C5 16'h806C
`define CUBE_LUT_A4C1 16'h806B
`define CUBE_LUT_A4BC 16'h806A
`define CUBE_LUT_A4B7 16'h8069
`define CUBE_LUT_A4B2 16'h8068
`define CUBE_LUT_A4AD 16'h8066
`define CUBE_LUT_A4A8 16'h8065
`define CUBE_LUT_A4A3 16'h8064
`define CUBE_LUT_A49E 16'h8062
`define CUBE_LUT_A499 16'h8061
`define CUBE_LUT_A494 16'h8060
`define CUBE_LUT_A48F 16'h805F
`define CUBE_LUT_A48A 16'h805E
`define CUBE_LUT_A486 16'h805D
`define CUBE_LUT_A481 16'h805B
`define CUBE_LUT_A47C 16'h805A
`define CUBE_LUT_A477 16'h8059
`define CUBE_LUT_A472 16'h8058
`define CUBE_LUT_A46D 16'h8057
`define CUBE_LUT_A468 16'h8056
`define CUBE_LUT_A463 16'h8054
`define CUBE_LUT_A45E 16'h8053
`define CUBE_LUT_A459 16'h8052
`define CUBE_LUT_A454 16'h8051
`define CUBE_LUT_A44F 16'h8050
`define CUBE_LUT_A44B 16'h804F
`define CUBE_LUT_A446 16'h804E
`define CUBE_LUT_A441 16'h804D
`define CUBE_LUT_A43C 16'h804C
`define CUBE_LUT_A437 16'h804B
`define CUBE_LUT_A432 16'h804A
`define CUBE_LUT_A42D 16'h8049
`define CUBE_LUT_A428 16'h8048
`define CUBE_LUT_A423 16'h8047
`define CUBE_LUT_A41E 16'h8046
`define CUBE_LUT_A419 16'h8045
`define CUBE_LUT_A414 16'h8044
`define CUBE_LUT_A410 16'h8043
`define CUBE_LUT_A40B 16'h8042
`define CUBE_LUT_A406 16'h8041
`define CUBE_LUT_A401 16'h8040
`define CUBE_LUT_A3F8 16'h803F
`define CUBE_LUT_A3EE 16'h803E
`define CUBE_LUT_A3E4 16'h803D
`define CUBE_LUT_A3DA 16'h803D
`define CUBE_LUT_A3D1 16'h803C
`define CUBE_LUT_A3C7 16'h803B
`define CUBE_LUT_A3BD 16'h803A
`define CUBE_LUT_A3B3 16'h8039
`define CUBE_LUT_A3A9 16'h8038
`define CUBE_LUT_A39F 16'h8037
`define CUBE_LUT_A396 16'h8037
`define CUBE_LUT_A38C 16'h8036
`define CUBE_LUT_A382 16'h8035
`define CUBE_LUT_A378 16'h8034
`define CUBE_LUT_A36E 16'h8033
`define CUBE_LUT_A364 16'h8032
`define CUBE_LUT_A35B 16'h8032
`define CUBE_LUT_A351 16'h8031
`define CUBE_LUT_A347 16'h8030
`define CUBE_LUT_A33D 16'h802F
`define CUBE_LUT_A333 16'h802F
`define CUBE_LUT_A329 16'h802E
`define CUBE_LUT_A320 16'h802D
`define CUBE_LUT_A316 16'h802C
`define CUBE_LUT_A30C 16'h802C
`define CUBE_LUT_A302 16'h802B
`define CUBE_LUT_A2F8 16'h802A
`define CUBE_LUT_A2EE 16'h802A
`define CUBE_LUT_A2E5 16'h8029
`define CUBE_LUT_A2DB 16'h8028
`define CUBE_LUT_A2D1 16'h8028
`define CUBE_LUT_A2C7 16'h8027
`define CUBE_LUT_A2BD 16'h8026
`define CUBE_LUT_A2B3 16'h8026
`define CUBE_LUT_A2AA 16'h8025
`define CUBE_LUT_A2A0 16'h8024
`define CUBE_LUT_A296 16'h8024
`define CUBE_LUT_A28C 16'h8023
`define CUBE_LUT_A282 16'h8022
`define CUBE_LUT_A278 16'h8022
`define CUBE_LUT_A26F 16'h8021
`define CUBE_LUT_A265 16'h8021
`define CUBE_LUT_A25B 16'h8020
`define CUBE_LUT_A251 16'h8020
`define CUBE_LUT_A247 16'h801F
`define CUBE_LUT_A23D 16'h801E
`define CUBE_LUT_A234 16'h801E
`define CUBE_LUT_A22A 16'h801D
`define CUBE_LUT_A220 16'h801D
`define CUBE_LUT_A216 16'h801C
`define CUBE_LUT_A20C 16'h801C
`define CUBE_LUT_A202 16'h801B
`define CUBE_LUT_A1F9 16'h801B
`define CUBE_LUT_A1EF 16'h801A
`define CUBE_LUT_A1E5 16'h801A
`define CUBE_LUT_A1DB 16'h8019
`define CUBE_LUT_A1D1 16'h8019
`define CUBE_LUT_A1C7 16'h8018
`define CUBE_LUT_A1BE 16'h8018
`define CUBE_LUT_A1B4 16'h8017
`define CUBE_LUT_A1AA 16'h8017
`define CUBE_LUT_A1A0 16'h8016
`define CUBE_LUT_A196 16'h8016
`define CUBE_LUT_A18D 16'h8015
`define CUBE_LUT_A183 16'h8015
`define CUBE_LUT_A179 16'h8014
`define CUBE_LUT_A16F 16'h8014
`define CUBE_LUT_A165 16'h8014
`define CUBE_LUT_A15B 16'h8013
`define CUBE_LUT_A152 16'h8013
`define CUBE_LUT_A148 16'h8012
`define CUBE_LUT_A13E 16'h8012
`define CUBE_LUT_A134 16'h8012
`define CUBE_LUT_A12A 16'h8011
`define CUBE_LUT_A120 16'h8011
`define CUBE_LUT_A117 16'h8010
`define CUBE_LUT_A10D 16'h8010
`define CUBE_LUT_A103 16'h8010
`define CUBE_LUT_A0F9 16'h800F
`define CUBE_LUT_A0EF 16'h800F
`define CUBE_LUT_A0E5 16'h800F
`define CUBE_LUT_A0DC 16'h800E
`define CUBE_LUT_A0D2 16'h800E
`define CUBE_LUT_A0C8 16'h800E
`define CUBE_LUT_A0BE 16'h800D
`define CUBE_LUT_A0B4 16'h800D
`define CUBE_LUT_A0AA 16'h800D
`define CUBE_LUT_A0A1 16'h800C
`define CUBE_LUT_A097 16'h800C
`define CUBE_LUT_A08D 16'h800C
`define CUBE_LUT_A083 16'h800B
`define CUBE_LUT_A079 16'h800B
`define CUBE_LUT_A06F 16'h800B
`define CUBE_LUT_A066 16'h800B
`define CUBE_LUT_A05C 16'h800A
`define CUBE_LUT_A052 16'h800A
`define CUBE_LUT_A048 16'h800A
`define CUBE_LUT_A03E 16'h800A
`define CUBE_LUT_A034 16'h8009
`define CUBE_LUT_A02B 16'h8009
`define CUBE_LUT_A021 16'h8009
`define CUBE_LUT_A017 16'h8009
`define CUBE_LUT_A00D 16'h8008
`define CUBE_LUT_A003 16'h8008
`define CUBE_LUT_9FF3 16'h8008
`define CUBE_LUT_9FDF 16'h8008
`define CUBE_LUT_9FCC 16'h8007
`define CUBE_LUT_9FB8 16'h8007
`define CUBE_LUT_9FA4 16'h8007
`define CUBE_LUT_9F91 16'h8007
`define CUBE_LUT_9F7D 16'h8007
`define CUBE_LUT_9F69 16'h8006
`define CUBE_LUT_9F56 16'h8006
`define CUBE_LUT_9F42 16'h8006
`define CUBE_LUT_9F2E 16'h8006
`define CUBE_LUT_9F1B 16'h8006
`define CUBE_LUT_9F07 16'h8005
`define CUBE_LUT_9EF3 16'h8005
`define CUBE_LUT_9EE0 16'h8005
`define CUBE_LUT_9ECC 16'h8005
`define CUBE_LUT_9EB8 16'h8005
`define CUBE_LUT_9EA5 16'h8005
`define CUBE_LUT_9E91 16'h8004
`define CUBE_LUT_9E7D 16'h8004
`define CUBE_LUT_9E6A 16'h8004
`define CUBE_LUT_9E56 16'h8004
`define CUBE_LUT_9E42 16'h8004
`define CUBE_LUT_9E2F 16'h8004
`define CUBE_LUT_9E1B 16'h8004
`define CUBE_LUT_9E07 16'h8003
`define CUBE_LUT_9DF4 16'h8003
`define CUBE_LUT_9DE0 16'h8003
`define CUBE_LUT_9DCC 16'h8003
`define CUBE_LUT_9DB9 16'h8003
`define CUBE_LUT_9DA5 16'h8003
`define CUBE_LUT_9D91 16'h8003
`define CUBE_LUT_9D7E 16'h8003
`define CUBE_LUT_9D6A 16'h8002
`define CUBE_LUT_9D56 16'h8002
`define CUBE_LUT_9D43 16'h8002
`define CUBE_LUT_9D2F 16'h8002
`define CUBE_LUT_9D1B 16'h8002
`define CUBE_LUT_9D08 16'h8002
`define CUBE_LUT_9CF4 16'h8002
`define CUBE_LUT_9CE0 16'h8002
`define CUBE_LUT_9CCD 16'h8002
`define CUBE_LUT_9CB9 16'h8002
`define CUBE_LUT_9CA5 16'h8002
`define CUBE_LUT_9C92 16'h8001
`define CUBE_LUT_9C7E 16'h8001
`define CUBE_LUT_9C6B 16'h8001
`define CUBE_LUT_9C57 16'h8001
`define CUBE_LUT_9C43 16'h8001
`define CUBE_LUT_9C30 16'h8001
`define CUBE_LUT_9C1C 16'h8001
`define CUBE_LUT_9C08 16'h8001
`define CUBE_LUT_9BE9 16'h8001
`define CUBE_LUT_9BC2 16'h8001
`define CUBE_LUT_9B9A 16'h8001
`define CUBE_LUT_9B73 16'h8001
`define CUBE_LUT_9B4C 16'h8001
`define CUBE_LUT_9B24 16'h8001
`define CUBE_LUT_9AFD 16'h8001
`define CUBE_LUT_9AD6 16'h8001
`define CUBE_LUT_9AAF 16'h8001
`define CUBE_LUT_9A87 16'h8001
`define CUBE_LUT_9A60 16'h8001
`define CUBE_LUT_9A39 16'h8000
`define CUBE_LUT_9A11 16'h8000
`define CUBE_LUT_99EA 16'h8000
`define CUBE_LUT_99C3 16'h8000
`define CUBE_LUT_999B 16'h8000
`define CUBE_LUT_9974 16'h8000
`define CUBE_LUT_994D 16'h8000
`define CUBE_LUT_9925 16'h8000
`define CUBE_LUT_98FE 16'h8000
`define CUBE_LUT_98D7 16'h8000
`define CUBE_LUT_98AF 16'h8000
`define CUBE_LUT_9888 16'h8000
`define CUBE_LUT_9861 16'h8000
`define CUBE_LUT_9839 16'h8000
`define CUBE_LUT_9812 16'h8000
`define CUBE_LUT_97D5 16'h8000
`define CUBE_LUT_9787 16'h8000
`define CUBE_LUT_9738 16'h8000
`define CUBE_LUT_96E9 16'h8000
`define CUBE_LUT_969B 16'h8000
`define CUBE_LUT_964C 16'h8000
`define CUBE_LUT_95FE 16'h8000
`define CUBE_LUT_95AF 16'h8000
`define CUBE_LUT_9560 16'h8000
`define CUBE_LUT_9512 16'h8000
`define CUBE_LUT_94C3 16'h8000
`define CUBE_LUT_9474 16'h8000
`define CUBE_LUT_9426 16'h8000
`define CUBE_LUT_93AE 16'h8000
`define CUBE_LUT_9311 16'h8000
`define CUBE_LUT_9274 16'h8000
`define CUBE_LUT_91D6 16'h8000
`define CUBE_LUT_9139 16'h8000
`define CUBE_LUT_909C 16'h8000
`define CUBE_LUT_8FFD 16'h8000
`define CUBE_LUT_8EC2 16'h8000
`define CUBE_LUT_8D88 16'h8000
`define CUBE_LUT_8C4D 16'h8000
`define CUBE_LUT_8A25 16'h8000
`define CUBE_LUT_875F 16'h8000
`define CUBE_LUT_8275 16'h8000
`define CUBE_LUT_0275 16'h0000
`define CUBE_LUT_075F 16'h0000
`define CUBE_LUT_0A25 16'h0000
`define CUBE_LUT_0C4D 16'h0000
`define CUBE_LUT_0D88 16'h0000
`define CUBE_LUT_0EC2 16'h0000
`define CUBE_LUT_0FFD 16'h0000
`define CUBE_LUT_109C 16'h0000
`define CUBE_LUT_1139 16'h0000
`define CUBE_LUT_11D6 16'h0000
`define CUBE_LUT_1274 16'h0000
`define CUBE_LUT_1311 16'h0000
`define CUBE_LUT_13AE 16'h0000
`define CUBE_LUT_1426 16'h0000
`define CUBE_LUT_1474 16'h0000
`define CUBE_LUT_14C3 16'h0000
`define CUBE_LUT_1512 16'h0000
`define CUBE_LUT_1560 16'h0000
`define CUBE_LUT_15AF 16'h0000
`define CUBE_LUT_15FE 16'h0000
`define CUBE_LUT_164C 16'h0000
`define CUBE_LUT_169B 16'h0000
`define CUBE_LUT_16E9 16'h0000
`define CUBE_LUT_1738 16'h0000
`define CUBE_LUT_1787 16'h0000
`define CUBE_LUT_17D5 16'h0000
`define CUBE_LUT_1812 16'h0000
`define CUBE_LUT_1839 16'h0000
`define CUBE_LUT_1861 16'h0000
`define CUBE_LUT_1888 16'h0000
`define CUBE_LUT_18AF 16'h0000
`define CUBE_LUT_18D7 16'h0000
`define CUBE_LUT_18FE 16'h0000
`define CUBE_LUT_1925 16'h0000
`define CUBE_LUT_194D 16'h0000
`define CUBE_LUT_1974 16'h0000
`define CUBE_LUT_199B 16'h0000
`define CUBE_LUT_19C3 16'h0000
`define CUBE_LUT_19EA 16'h0000
`define CUBE_LUT_1A11 16'h0000
`define CUBE_LUT_1A39 16'h0000
`define CUBE_LUT_1A60 16'h0001
`define CUBE_LUT_1A87 16'h0001
`define CUBE_LUT_1AAF 16'h0001
`define CUBE_LUT_1AD6 16'h0001
`define CUBE_LUT_1AFD 16'h0001
`define CUBE_LUT_1B24 16'h0001
`define CUBE_LUT_1B4C 16'h0001
`define CUBE_LUT_1B73 16'h0001
`define CUBE_LUT_1B9A 16'h0001
`define CUBE_LUT_1BC2 16'h0001
`define CUBE_LUT_1BE9 16'h0001
`define CUBE_LUT_1C08 16'h0001
`define CUBE_LUT_1C1C 16'h0001
`define CUBE_LUT_1C30 16'h0001
`define CUBE_LUT_1C43 16'h0001
`define CUBE_LUT_1C57 16'h0001
`define CUBE_LUT_1C6B 16'h0001
`define CUBE_LUT_1C7E 16'h0001
`define CUBE_LUT_1C92 16'h0001
`define CUBE_LUT_1CA5 16'h0002
`define CUBE_LUT_1CB9 16'h0002
`define CUBE_LUT_1CCD 16'h0002
`define CUBE_LUT_1CE0 16'h0002
`define CUBE_LUT_1CF4 16'h0002
`define CUBE_LUT_1D08 16'h0002
`define CUBE_LUT_1D1B 16'h0002
`define CUBE_LUT_1D2F 16'h0002
`define CUBE_LUT_1D43 16'h0002
`define CUBE_LUT_1D56 16'h0002
`define CUBE_LUT_1D6A 16'h0002
`define CUBE_LUT_1D7E 16'h0003
`define CUBE_LUT_1D91 16'h0003
`define CUBE_LUT_1DA5 16'h0003
`define CUBE_LUT_1DB9 16'h0003
`define CUBE_LUT_1DCC 16'h0003
`define CUBE_LUT_1DE0 16'h0003
`define CUBE_LUT_1DF4 16'h0003
`define CUBE_LUT_1E07 16'h0003
`define CUBE_LUT_1E1B 16'h0004
`define CUBE_LUT_1E2F 16'h0004
`define CUBE_LUT_1E42 16'h0004
`define CUBE_LUT_1E56 16'h0004
`define CUBE_LUT_1E6A 16'h0004
`define CUBE_LUT_1E7D 16'h0004
`define CUBE_LUT_1E91 16'h0004
`define CUBE_LUT_1EA5 16'h0005
`define CUBE_LUT_1EB8 16'h0005
`define CUBE_LUT_1ECC 16'h0005
`define CUBE_LUT_1EE0 16'h0005
`define CUBE_LUT_1EF3 16'h0005
`define CUBE_LUT_1F07 16'h0005
`define CUBE_LUT_1F1B 16'h0006
`define CUBE_LUT_1F2E 16'h0006
`define CUBE_LUT_1F42 16'h0006
`define CUBE_LUT_1F56 16'h0006
`define CUBE_LUT_1F69 16'h0006
`define CUBE_LUT_1F7D 16'h0007
`define CUBE_LUT_1F91 16'h0007
`define CUBE_LUT_1FA4 16'h0007
`define CUBE_LUT_1FB8 16'h0007
`define CUBE_LUT_1FCC 16'h0007
`define CUBE_LUT_1FDF 16'h0008
`define CUBE_LUT_1FF3 16'h0008
`define CUBE_LUT_2003 16'h0008
`define CUBE_LUT_200D 16'h0008
`define CUBE_LUT_2017 16'h0009
`define CUBE_LUT_2021 16'h0009
`define CUBE_LUT_202B 16'h0009
`define CUBE_LUT_2034 16'h0009
`define CUBE_LUT_203E 16'h000A
`define CUBE_LUT_2048 16'h000A
`define CUBE_LUT_2052 16'h000A
`define CUBE_LUT_205C 16'h000A
`define CUBE_LUT_2066 16'h000B
`define CUBE_LUT_206F 16'h000B
`define CUBE_LUT_2079 16'h000B
`define CUBE_LUT_2083 16'h000B
`define CUBE_LUT_208D 16'h000C
`define CUBE_LUT_2097 16'h000C
`define CUBE_LUT_20A1 16'h000C
`define CUBE_LUT_20AA 16'h000D
`define CUBE_LUT_20B4 16'h000D
`define CUBE_LUT_20BE 16'h000D
`define CUBE_LUT_20C8 16'h000E
`define CUBE_LUT_20D2 16'h000E
`define CUBE_LUT_20DC 16'h000E
`define CUBE_LUT_20E5 16'h000F
`define CUBE_LUT_20EF 16'h000F
`define CUBE_LUT_20F9 16'h000F
`define CUBE_LUT_2103 16'h0010
`define CUBE_LUT_210D 16'h0010
`define CUBE_LUT_2117 16'h0010
`define CUBE_LUT_2120 16'h0011
`define CUBE_LUT_212A 16'h0011
`define CUBE_LUT_2134 16'h0012
`define CUBE_LUT_213E 16'h0012
`define CUBE_LUT_2148 16'h0012
`define CUBE_LUT_2152 16'h0013
`define CUBE_LUT_215B 16'h0013
`define CUBE_LUT_2165 16'h0014
`define CUBE_LUT_216F 16'h0014
`define CUBE_LUT_2179 16'h0014
`define CUBE_LUT_2183 16'h0015
`define CUBE_LUT_218D 16'h0015
`define CUBE_LUT_2196 16'h0016
`define CUBE_LUT_21A0 16'h0016
`define CUBE_LUT_21AA 16'h0017
`define CUBE_LUT_21B4 16'h0017
`define CUBE_LUT_21BE 16'h0018
`define CUBE_LUT_21C7 16'h0018
`define CUBE_LUT_21D1 16'h0019
`define CUBE_LUT_21DB 16'h0019
`define CUBE_LUT_21E5 16'h001A
`define CUBE_LUT_21EF 16'h001A
`define CUBE_LUT_21F9 16'h001B
`define CUBE_LUT_2202 16'h001B
`define CUBE_LUT_220C 16'h001C
`define CUBE_LUT_2216 16'h001C
`define CUBE_LUT_2220 16'h001D
`define CUBE_LUT_222A 16'h001D
`define CUBE_LUT_2234 16'h001E
`define CUBE_LUT_223D 16'h001E
`define CUBE_LUT_2247 16'h001F
`define CUBE_LUT_2251 16'h0020
`define CUBE_LUT_225B 16'h0020
`define CUBE_LUT_2265 16'h0021
`define CUBE_LUT_226F 16'h0021
`define CUBE_LUT_2278 16'h0022
`define CUBE_LUT_2282 16'h0022
`define CUBE_LUT_228C 16'h0023
`define CUBE_LUT_2296 16'h0024
`define CUBE_LUT_22A0 16'h0024
`define CUBE_LUT_22AA 16'h0025
`define CUBE_LUT_22B3 16'h0026
`define CUBE_LUT_22BD 16'h0026
`define CUBE_LUT_22C7 16'h0027
`define CUBE_LUT_22D1 16'h0028
`define CUBE_LUT_22DB 16'h0028
`define CUBE_LUT_22E5 16'h0029
`define CUBE_LUT_22EE 16'h002A
`define CUBE_LUT_22F8 16'h002A
`define CUBE_LUT_2302 16'h002B
`define CUBE_LUT_230C 16'h002C
`define CUBE_LUT_2316 16'h002C
`define CUBE_LUT_2320 16'h002D
`define CUBE_LUT_2329 16'h002E
`define CUBE_LUT_2333 16'h002F
`define CUBE_LUT_233D 16'h002F
`define CUBE_LUT_2347 16'h0030
`define CUBE_LUT_2351 16'h0031
`define CUBE_LUT_235B 16'h0032
`define CUBE_LUT_2364 16'h0032
`define CUBE_LUT_236E 16'h0033
`define CUBE_LUT_2378 16'h0034
`define CUBE_LUT_2382 16'h0035
`define CUBE_LUT_238C 16'h0036
`define CUBE_LUT_2396 16'h0037
`define CUBE_LUT_239F 16'h0037
`define CUBE_LUT_23A9 16'h0038
`define CUBE_LUT_23B3 16'h0039
`define CUBE_LUT_23BD 16'h003A
`define CUBE_LUT_23C7 16'h003B
`define CUBE_LUT_23D1 16'h003C
`define CUBE_LUT_23DA 16'h003D
`define CUBE_LUT_23E4 16'h003D
`define CUBE_LUT_23EE 16'h003E
`define CUBE_LUT_23F8 16'h003F
`define CUBE_LUT_2401 16'h0040
`define CUBE_LUT_2406 16'h0041
`define CUBE_LUT_240B 16'h0042
`define CUBE_LUT_2410 16'h0043
`define CUBE_LUT_2414 16'h0044
`define CUBE_LUT_2419 16'h0045
`define CUBE_LUT_241E 16'h0046
`define CUBE_LUT_2423 16'h0047
`define CUBE_LUT_2428 16'h0048
`define CUBE_LUT_242D 16'h0049
`define CUBE_LUT_2432 16'h004A
`define CUBE_LUT_2437 16'h004B
`define CUBE_LUT_243C 16'h004C
`define CUBE_LUT_2441 16'h004D
`define CUBE_LUT_2446 16'h004E
`define CUBE_LUT_244B 16'h004F
`define CUBE_LUT_244F 16'h0050
`define CUBE_LUT_2454 16'h0051
`define CUBE_LUT_2459 16'h0052
`define CUBE_LUT_245E 16'h0053
`define CUBE_LUT_2463 16'h0054
`define CUBE_LUT_2468 16'h0056
`define CUBE_LUT_246D 16'h0057
`define CUBE_LUT_2472 16'h0058
`define CUBE_LUT_2477 16'h0059
`define CUBE_LUT_247C 16'h005A
`define CUBE_LUT_2481 16'h005B
`define CUBE_LUT_2486 16'h005D
`define CUBE_LUT_248A 16'h005E
`define CUBE_LUT_248F 16'h005F
`define CUBE_LUT_2494 16'h0060
`define CUBE_LUT_2499 16'h0061
`define CUBE_LUT_249E 16'h0062
`define CUBE_LUT_24A3 16'h0064
`define CUBE_LUT_24A8 16'h0065
`define CUBE_LUT_24AD 16'h0066
`define CUBE_LUT_24B2 16'h0068
`define CUBE_LUT_24B7 16'h0069
`define CUBE_LUT_24BC 16'h006A
`define CUBE_LUT_24C1 16'h006B
`define CUBE_LUT_24C5 16'h006C
`define CUBE_LUT_24CA 16'h006E
`define CUBE_LUT_24CF 16'h006F
`define CUBE_LUT_24D4 16'h0071
`define CUBE_LUT_24D9 16'h0072
`define CUBE_LUT_24DE 16'h0073
`define CUBE_LUT_24E3 16'h0075
`define CUBE_LUT_24E8 16'h0076
`define CUBE_LUT_24ED 16'h0078
`define CUBE_LUT_24F2 16'h0079
`define CUBE_LUT_24F7 16'h007A
`define CUBE_LUT_24FC 16'h007C
`define CUBE_LUT_2500 16'h007D
`define CUBE_LUT_2505 16'h007E
`define CUBE_LUT_250A 16'h0080
`define CUBE_LUT_250F 16'h0081
`define CUBE_LUT_2514 16'h0083
`define CUBE_LUT_2519 16'h0084
`define CUBE_LUT_251E 16'h0086
`define CUBE_LUT_2523 16'h0088
`define CUBE_LUT_2528 16'h0089
`define CUBE_LUT_252D 16'h008B
`define CUBE_LUT_2532 16'h008C
`define CUBE_LUT_2536 16'h008D
`define CUBE_LUT_253B 16'h008F
`define CUBE_LUT_2540 16'h0091
`define CUBE_LUT_2545 16'h0092
`define CUBE_LUT_254A 16'h0094
`define CUBE_LUT_254F 16'h0096
`define CUBE_LUT_2554 16'h0097
`define CUBE_LUT_2559 16'h0099
`define CUBE_LUT_255E 16'h009B
`define CUBE_LUT_2563 16'h009C
`define CUBE_LUT_2568 16'h009E
`define CUBE_LUT_256D 16'h00A0
`define CUBE_LUT_2571 16'h00A1
`define CUBE_LUT_2576 16'h00A3
`define CUBE_LUT_257B 16'h00A5
`define CUBE_LUT_2580 16'h00A6
`define CUBE_LUT_2585 16'h00A8
`define CUBE_LUT_258A 16'h00AA
`define CUBE_LUT_258F 16'h00AC
`define CUBE_LUT_2594 16'h00AE
`define CUBE_LUT_2599 16'h00AF
`define CUBE_LUT_259E 16'h00B1
`define CUBE_LUT_25A3 16'h00B3
`define CUBE_LUT_25A8 16'h00B5
`define CUBE_LUT_25AC 16'h00B6
`define CUBE_LUT_25B1 16'h00B8
`define CUBE_LUT_25B6 16'h00BA
`define CUBE_LUT_25BB 16'h00BC
`define CUBE_LUT_25C0 16'h00BE
`define CUBE_LUT_25C5 16'h00C0
`define CUBE_LUT_25CA 16'h00C2
`define CUBE_LUT_25CF 16'h00C4
`define CUBE_LUT_25D4 16'h00C6
`define CUBE_LUT_25D9 16'h00C8
`define CUBE_LUT_25DE 16'h00CA
`define CUBE_LUT_25E3 16'h00CC
`define CUBE_LUT_25E7 16'h00CE
`define CUBE_LUT_25EC 16'h00D0
`define CUBE_LUT_25F1 16'h00D2
`define CUBE_LUT_25F6 16'h00D4
`define CUBE_LUT_25FB 16'h00D6
`define CUBE_LUT_2600 16'h00D8
`define CUBE_LUT_2605 16'h00DA
`define CUBE_LUT_260A 16'h00DC
`define CUBE_LUT_260F 16'h00DE
`define CUBE_LUT_2614 16'h00E1
`define CUBE_LUT_2619 16'h00E3
`define CUBE_LUT_261E 16'h00E5
`define CUBE_LUT_2622 16'h00E7
`define CUBE_LUT_2627 16'h00E9
`define CUBE_LUT_262C 16'h00EB
`define CUBE_LUT_2631 16'h00ED
`define CUBE_LUT_2636 16'h00F0
`define CUBE_LUT_263B 16'h00F2
`define CUBE_LUT_2640 16'h00F4
`define CUBE_LUT_2645 16'h00F6
`define CUBE_LUT_264A 16'h00F9
`define CUBE_LUT_264F 16'h00FB
`define CUBE_LUT_2654 16'h00FD
`define CUBE_LUT_2658 16'h00FF
`define CUBE_LUT_265D 16'h0102
`define CUBE_LUT_2662 16'h0104
`define CUBE_LUT_2667 16'h0106
`define CUBE_LUT_266C 16'h0109
`define CUBE_LUT_2671 16'h010B
`define CUBE_LUT_2676 16'h010E
`define CUBE_LUT_267B 16'h0110
`define CUBE_LUT_2680 16'h0113
`define CUBE_LUT_2685 16'h0115
`define CUBE_LUT_268A 16'h0118
`define CUBE_LUT_268F 16'h011A
`define CUBE_LUT_2693 16'h011C
`define CUBE_LUT_2698 16'h011F
`define CUBE_LUT_269D 16'h0121
`define CUBE_LUT_26A2 16'h0124
`define CUBE_LUT_26A7 16'h0126
`define CUBE_LUT_26AC 16'h0129
`define CUBE_LUT_26B1 16'h012C
`define CUBE_LUT_26B6 16'h012E
`define CUBE_LUT_26BB 16'h0131
`define CUBE_LUT_26C0 16'h0134
`define CUBE_LUT_26C5 16'h0136
`define CUBE_LUT_26CA 16'h0139
`define CUBE_LUT_26CE 16'h013B
`define CUBE_LUT_26D3 16'h013E
`define CUBE_LUT_26D8 16'h0141
`define CUBE_LUT_26DD 16'h0143
`define CUBE_LUT_26E2 16'h0146
`define CUBE_LUT_26E7 16'h0149
`define CUBE_LUT_26EC 16'h014C
`define CUBE_LUT_26F1 16'h014E
`define CUBE_LUT_26F6 16'h0151
`define CUBE_LUT_26FB 16'h0154
`define CUBE_LUT_2700 16'h0157
`define CUBE_LUT_2705 16'h015A
`define CUBE_LUT_2709 16'h015C
`define CUBE_LUT_270E 16'h015F
`define CUBE_LUT_2713 16'h0162
`define CUBE_LUT_2718 16'h0165
`define CUBE_LUT_271D 16'h0168
`define CUBE_LUT_2722 16'h016B
`define CUBE_LUT_2727 16'h016E
`define CUBE_LUT_272C 16'h0171
`define CUBE_LUT_2731 16'h0174
`define CUBE_LUT_2736 16'h0177
`define CUBE_LUT_273B 16'h017A
`define CUBE_LUT_2740 16'h017D
`define CUBE_LUT_2744 16'h0180
`define CUBE_LUT_2749 16'h0183
`define CUBE_LUT_274E 16'h0186
`define CUBE_LUT_2753 16'h0189
`define CUBE_LUT_2758 16'h018C
`define CUBE_LUT_275D 16'h018F
`define CUBE_LUT_2762 16'h0192
`define CUBE_LUT_2767 16'h0196
`define CUBE_LUT_276C 16'h0199
`define CUBE_LUT_2771 16'h019C
`define CUBE_LUT_2776 16'h019F
`define CUBE_LUT_277A 16'h01A2
`define CUBE_LUT_277F 16'h01A5
`define CUBE_LUT_2784 16'h01A9
`define CUBE_LUT_2789 16'h01AC
`define CUBE_LUT_278E 16'h01AF
`define CUBE_LUT_2793 16'h01B3
`define CUBE_LUT_2798 16'h01B6
`define CUBE_LUT_279D 16'h01B9
`define CUBE_LUT_27A2 16'h01BD
`define CUBE_LUT_27A7 16'h01C0
`define CUBE_LUT_27AC 16'h01C4
`define CUBE_LUT_27B1 16'h01C7
`define CUBE_LUT_27B5 16'h01CA
`define CUBE_LUT_27BA 16'h01CD
`define CUBE_LUT_27BF 16'h01D1
`define CUBE_LUT_27C4 16'h01D4
`define CUBE_LUT_27C9 16'h01D8
`define CUBE_LUT_27CE 16'h01DB
`define CUBE_LUT_27D3 16'h01DF
`define CUBE_LUT_27D8 16'h01E3
`define CUBE_LUT_27DD 16'h01E6
`define CUBE_LUT_27E2 16'h01EA
`define CUBE_LUT_27E7 16'h01ED
`define CUBE_LUT_27EC 16'h01F1
`define CUBE_LUT_27F0 16'h01F4
`define CUBE_LUT_27F5 16'h01F8
`define CUBE_LUT_27FA 16'h01FC
`define CUBE_LUT_27FF 16'h01FF
`define CUBE_LUT_2802 16'h0203
`define CUBE_LUT_2805 16'h0208
`define CUBE_LUT_2807 16'h020B
`define CUBE_LUT_2809 16'h020E
`define CUBE_LUT_280C 16'h0212
`define CUBE_LUT_280E 16'h0215
`define CUBE_LUT_2811 16'h021A
`define CUBE_LUT_2813 16'h021D
`define CUBE_LUT_2816 16'h0222
`define CUBE_LUT_2818 16'h0225
`define CUBE_LUT_281B 16'h022A
`define CUBE_LUT_281D 16'h022D
`define CUBE_LUT_2820 16'h0232
`define CUBE_LUT_2822 16'h0235
`define CUBE_LUT_2824 16'h0238
`define CUBE_LUT_2827 16'h023D
`define CUBE_LUT_2829 16'h0240
`define CUBE_LUT_282C 16'h0245
`define CUBE_LUT_282E 16'h0248
`define CUBE_LUT_2831 16'h024D
`define CUBE_LUT_2833 16'h0250
`define CUBE_LUT_2836 16'h0255
`define CUBE_LUT_2838 16'h0259
`define CUBE_LUT_283B 16'h025E
`define CUBE_LUT_283D 16'h0261
`define CUBE_LUT_2840 16'h0266
`define CUBE_LUT_2842 16'h026A
`define CUBE_LUT_2844 16'h026D
`define CUBE_LUT_2847 16'h0272
`define CUBE_LUT_2849 16'h0275
`define CUBE_LUT_284C 16'h027B
`define CUBE_LUT_284E 16'h027E
`define CUBE_LUT_2851 16'h0283
`define CUBE_LUT_2853 16'h0287
`define CUBE_LUT_2856 16'h028C
`define CUBE_LUT_2858 16'h0290
`define CUBE_LUT_285B 16'h0295
`define CUBE_LUT_285D 16'h0299
`define CUBE_LUT_285F 16'h029C
`define CUBE_LUT_2862 16'h02A2
`define CUBE_LUT_2864 16'h02A5
`define CUBE_LUT_2867 16'h02AB
`define CUBE_LUT_2869 16'h02AE
`define CUBE_LUT_286C 16'h02B4
`define CUBE_LUT_286E 16'h02B7
`define CUBE_LUT_2871 16'h02BD
`define CUBE_LUT_2873 16'h02C1
`define CUBE_LUT_2876 16'h02C6
`define CUBE_LUT_2878 16'h02CA
`define CUBE_LUT_287A 16'h02CE
`define CUBE_LUT_287D 16'h02D3
`define CUBE_LUT_287F 16'h02D7
`define CUBE_LUT_2882 16'h02DD
`define CUBE_LUT_2884 16'h02E1
`define CUBE_LUT_2887 16'h02E6
`define CUBE_LUT_2889 16'h02EA
`define CUBE_LUT_288C 16'h02F0
`define CUBE_LUT_288E 16'h02F4
`define CUBE_LUT_2891 16'h02FA
`define CUBE_LUT_2893 16'h02FE
`define CUBE_LUT_2896 16'h0304
`define CUBE_LUT_2898 16'h0308
`define CUBE_LUT_289A 16'h030B
`define CUBE_LUT_289D 16'h0311
`define CUBE_LUT_289F 16'h0315
`define CUBE_LUT_28A2 16'h031B
`define CUBE_LUT_28A4 16'h0320
`define CUBE_LUT_28A7 16'h0326
`define CUBE_LUT_28A9 16'h032A
`define CUBE_LUT_28AC 16'h0330
`define CUBE_LUT_28AE 16'h0334
`define CUBE_LUT_28B1 16'h033A
`define CUBE_LUT_28B3 16'h033E
`define CUBE_LUT_28B5 16'h0342
`define CUBE_LUT_28B8 16'h0349
`define CUBE_LUT_28BA 16'h034D
`define CUBE_LUT_28BD 16'h0353
`define CUBE_LUT_28BF 16'h0357
`define CUBE_LUT_28C2 16'h035E
`define CUBE_LUT_28C4 16'h0362
`define CUBE_LUT_28C7 16'h0368
`define CUBE_LUT_28C9 16'h036D
`define CUBE_LUT_28CC 16'h0373
`define CUBE_LUT_28CE 16'h0377
`define CUBE_LUT_28D1 16'h037E
`define CUBE_LUT_28D3 16'h0382
`define CUBE_LUT_28D5 16'h0387
`define CUBE_LUT_28D8 16'h038D
`define CUBE_LUT_28DA 16'h0392
`define CUBE_LUT_28DD 16'h0398
`define CUBE_LUT_28DF 16'h039D
`define CUBE_LUT_28E2 16'h03A3
`define CUBE_LUT_28E4 16'h03A8
`define CUBE_LUT_28E7 16'h03AF
`define CUBE_LUT_28E9 16'h03B3
`define CUBE_LUT_28EC 16'h03BA
`define CUBE_LUT_28EE 16'h03BE
`define CUBE_LUT_28F0 16'h03C3
`define CUBE_LUT_28F3 16'h03CA
`define CUBE_LUT_28F5 16'h03CE
`define CUBE_LUT_28F8 16'h03D5
`define CUBE_LUT_28FA 16'h03DA
`define CUBE_LUT_28FD 16'h03E1
`define CUBE_LUT_28FF 16'h03E6
`define CUBE_LUT_2902 16'h03ED
`define CUBE_LUT_2904 16'h03F1
`define CUBE_LUT_2907 16'h03F8
`define CUBE_LUT_2909 16'h03FD
`define CUBE_LUT_290B 16'h0402
`define CUBE_LUT_290E 16'h0409
`define CUBE_LUT_2910 16'h040E
`define CUBE_LUT_2913 16'h0415
`define CUBE_LUT_2915 16'h041A
`define CUBE_LUT_2918 16'h0421
`define CUBE_LUT_291A 16'h0426
`define CUBE_LUT_291D 16'h042E
`define CUBE_LUT_291F 16'h0432
`define CUBE_LUT_2922 16'h043A
`define CUBE_LUT_2924 16'h043F
`define CUBE_LUT_2927 16'h0446
`define CUBE_LUT_2929 16'h044B
`define CUBE_LUT_292B 16'h0450
`define CUBE_LUT_292E 16'h0458
`define CUBE_LUT_2930 16'h045D
`define CUBE_LUT_2933 16'h0464
`define CUBE_LUT_2935 16'h0469
`define CUBE_LUT_2938 16'h0471
`define CUBE_LUT_293A 16'h0476
`define CUBE_LUT_293D 16'h047E
`define CUBE_LUT_293F 16'h0483
`define CUBE_LUT_2942 16'h048B
`define CUBE_LUT_2944 16'h0490
`define CUBE_LUT_2946 16'h0495
`define CUBE_LUT_2949 16'h049D
`define CUBE_LUT_294B 16'h04A2
`define CUBE_LUT_294E 16'h04AA
`define CUBE_LUT_2950 16'h04AF
`define CUBE_LUT_2953 16'h04B7
`define CUBE_LUT_2955 16'h04BD
`define CUBE_LUT_2958 16'h04C5
`define CUBE_LUT_295A 16'h04CA
`define CUBE_LUT_295D 16'h04D2
`define CUBE_LUT_295F 16'h04D8
`define CUBE_LUT_2962 16'h04E0
`define CUBE_LUT_2964 16'h04E5
`define CUBE_LUT_2966 16'h04EB
`define CUBE_LUT_2969 16'h04F3
`define CUBE_LUT_296B 16'h04F8
`define CUBE_LUT_296E 16'h0501
`define CUBE_LUT_2970 16'h0506
`define CUBE_LUT_2973 16'h050E
`define CUBE_LUT_2975 16'h0514
`define CUBE_LUT_2978 16'h051C
`define CUBE_LUT_297A 16'h0522
`define CUBE_LUT_297D 16'h052B
`define CUBE_LUT_297F 16'h0530
`define CUBE_LUT_2981 16'h0536
`define CUBE_LUT_2984 16'h053E
`define CUBE_LUT_2986 16'h0544
`define CUBE_LUT_2989 16'h054D
`define CUBE_LUT_298B 16'h0552
`define CUBE_LUT_298E 16'h055B
`define CUBE_LUT_2990 16'h0561
`define CUBE_LUT_2993 16'h056A
`define CUBE_LUT_2995 16'h056F
`define CUBE_LUT_2998 16'h0578
`define CUBE_LUT_299A 16'h057E
`define CUBE_LUT_299C 16'h0584
`define CUBE_LUT_299F 16'h058D
`define CUBE_LUT_29A1 16'h0593
`define CUBE_LUT_29A4 16'h059C
`define CUBE_LUT_29A6 16'h05A2
`define CUBE_LUT_29A9 16'h05AB
`define CUBE_LUT_29AB 16'h05B1
`define CUBE_LUT_29AE 16'h05BA
`define CUBE_LUT_29B0 16'h05C0
`define CUBE_LUT_29B3 16'h05C9
`define CUBE_LUT_29B5 16'h05CF
`define CUBE_LUT_29B8 16'h05D8
`define CUBE_LUT_29BA 16'h05DE
`define CUBE_LUT_29BC 16'h05E5
`define CUBE_LUT_29BF 16'h05EE
`define CUBE_LUT_29C1 16'h05F4
`define CUBE_LUT_29C4 16'h05FD
`define CUBE_LUT_29C6 16'h0604
`define CUBE_LUT_29C9 16'h060D
`define CUBE_LUT_29CB 16'h0613
`define CUBE_LUT_29CE 16'h061D
`define CUBE_LUT_29D0 16'h0623
`define CUBE_LUT_29D3 16'h062D
`define CUBE_LUT_29D5 16'h0633
`define CUBE_LUT_29D7 16'h0639
`define CUBE_LUT_29DA 16'h0643
`define CUBE_LUT_29DC 16'h0649
`define CUBE_LUT_29DF 16'h0653
`define CUBE_LUT_29E1 16'h0659
`define CUBE_LUT_29E4 16'h0663
`define CUBE_LUT_29E6 16'h066A
`define CUBE_LUT_29E9 16'h0674
`define CUBE_LUT_29EB 16'h067A
`define CUBE_LUT_29EE 16'h0684
`define CUBE_LUT_29F0 16'h068B
`define CUBE_LUT_29F3 16'h0694
`define CUBE_LUT_29F5 16'h069B
`define CUBE_LUT_29F7 16'h06A2
`define CUBE_LUT_29FA 16'h06AC
`define CUBE_LUT_29FC 16'h06B3
`define CUBE_LUT_29FF 16'h06BD
`define CUBE_LUT_2A01 16'h06C3
`define CUBE_LUT_2A04 16'h06CE
`define CUBE_LUT_2A06 16'h06D4
`define CUBE_LUT_2A09 16'h06DF
`define CUBE_LUT_2A0B 16'h06E5
`define CUBE_LUT_2A0E 16'h06F0
`define CUBE_LUT_2A10 16'h06F7
`define CUBE_LUT_2A12 16'h06FD
`define CUBE_LUT_2A15 16'h0708
`define CUBE_LUT_2A17 16'h070F
`define CUBE_LUT_2A1A 16'h0719
`define CUBE_LUT_2A1C 16'h0720
`define CUBE_LUT_2A1F 16'h072B
`define CUBE_LUT_2A21 16'h0732
`define CUBE_LUT_2A24 16'h073C
`define CUBE_LUT_2A26 16'h0743
`define CUBE_LUT_2A29 16'h074E
`define CUBE_LUT_2A2B 16'h0755
`define CUBE_LUT_2A2D 16'h075C
`define CUBE_LUT_2A30 16'h0767
`define CUBE_LUT_2A32 16'h076E
`define CUBE_LUT_2A35 16'h0779
`define CUBE_LUT_2A37 16'h0780
`define CUBE_LUT_2A3A 16'h078B
`define CUBE_LUT_2A3C 16'h0793
`define CUBE_LUT_2A3F 16'h079D
`define CUBE_LUT_2A41 16'h07A5
`define CUBE_LUT_2A44 16'h07B0
`define CUBE_LUT_2A46 16'h07B7
`define CUBE_LUT_2A49 16'h07C2
`define CUBE_LUT_2A4B 16'h07CA
`define CUBE_LUT_2A4D 16'h07D1
`define CUBE_LUT_2A50 16'h07DC
`define CUBE_LUT_2A52 16'h07E4
`define CUBE_LUT_2A55 16'h07EF
`define CUBE_LUT_2A57 16'h07F7
`define CUBE_LUT_2A5A 16'h0801
`define CUBE_LUT_2A5C 16'h0805
`define CUBE_LUT_2A5F 16'h080A
`define CUBE_LUT_2A61 16'h080E
`define CUBE_LUT_2A64 16'h0814
`define CUBE_LUT_2A66 16'h0818
`define CUBE_LUT_2A68 16'h081C
`define CUBE_LUT_2A6B 16'h0821
`define CUBE_LUT_2A6D 16'h0825
`define CUBE_LUT_2A70 16'h082B
`define CUBE_LUT_2A72 16'h082F
`define CUBE_LUT_2A75 16'h0835
`define CUBE_LUT_2A77 16'h0839
`define CUBE_LUT_2A7A 16'h083F
`define CUBE_LUT_2A7C 16'h0843
`define CUBE_LUT_2A7F 16'h0849
`define CUBE_LUT_2A81 16'h084C
`define CUBE_LUT_2A84 16'h0852
`define CUBE_LUT_2A86 16'h0856
`define CUBE_LUT_2A88 16'h085A
`define CUBE_LUT_2A8B 16'h0860
`define CUBE_LUT_2A8D 16'h0864
`define CUBE_LUT_2A90 16'h086A
`define CUBE_LUT_2A92 16'h086F
`define CUBE_LUT_2A95 16'h0875
`define CUBE_LUT_2A97 16'h0879
`define CUBE_LUT_2A9A 16'h087F
`define CUBE_LUT_2A9C 16'h0883
`define CUBE_LUT_2A9F 16'h0889
`define CUBE_LUT_2AA1 16'h088D
`define CUBE_LUT_2AA3 16'h0891
`define CUBE_LUT_2AA6 16'h0897
`define CUBE_LUT_2AA8 16'h089C
`define CUBE_LUT_2AAB 16'h08A2
`define CUBE_LUT_2AAD 16'h08A6
`define CUBE_LUT_2AB0 16'h08AC
`define CUBE_LUT_2AB2 16'h08B1
`define CUBE_LUT_2AB5 16'h08B7
`define CUBE_LUT_2AB7 16'h08BB
`define CUBE_LUT_2ABA 16'h08C1
`define CUBE_LUT_2ABC 16'h08C6
`define CUBE_LUT_2ABE 16'h08CA
`define CUBE_LUT_2AC1 16'h08D0
`define CUBE_LUT_2AC3 16'h08D5
`define CUBE_LUT_2AC6 16'h08DB
`define CUBE_LUT_2AC8 16'h08DF
`define CUBE_LUT_2ACB 16'h08E6
`define CUBE_LUT_2ACD 16'h08EA
`define CUBE_LUT_2AD0 16'h08F1
`define CUBE_LUT_2AD2 16'h08F5
`define CUBE_LUT_2AD5 16'h08FC
`define CUBE_LUT_2AD7 16'h0900
`define CUBE_LUT_2ADA 16'h0907
`define CUBE_LUT_2ADC 16'h090B
`define CUBE_LUT_2ADE 16'h090F
`define CUBE_LUT_2AE1 16'h0916
`define CUBE_LUT_2AE3 16'h091A
`define CUBE_LUT_2AE6 16'h0921
`define CUBE_LUT_2AE8 16'h0926
`define CUBE_LUT_2AEB 16'h092C
`define CUBE_LUT_2AED 16'h0931
`define CUBE_LUT_2AF0 16'h0938
`define CUBE_LUT_2AF2 16'h093C
`define CUBE_LUT_2AF5 16'h0943
`define CUBE_LUT_2AF7 16'h0947
`define CUBE_LUT_2AF9 16'h094C
`define CUBE_LUT_2AFC 16'h0953
`define CUBE_LUT_2AFE 16'h0957
`define CUBE_LUT_2B01 16'h095E
`define CUBE_LUT_2B03 16'h0963
`define CUBE_LUT_2B06 16'h096A
`define CUBE_LUT_2B08 16'h096E
`define CUBE_LUT_2B0B 16'h0975
`define CUBE_LUT_2B0D 16'h097A
`define CUBE_LUT_2B10 16'h0981
`define CUBE_LUT_2B12 16'h0986
`define CUBE_LUT_2B15 16'h098D
`define CUBE_LUT_2B17 16'h0992
`define CUBE_LUT_2B19 16'h0996
`define CUBE_LUT_2B1C 16'h099D
`define CUBE_LUT_2B1E 16'h09A2
`define CUBE_LUT_2B21 16'h09A9
`define CUBE_LUT_2B23 16'h09AE
`define CUBE_LUT_2B26 16'h09B5
`define CUBE_LUT_2B28 16'h09BA
`define CUBE_LUT_2B2B 16'h09C1
`define CUBE_LUT_2B2D 16'h09C6
`define CUBE_LUT_2B30 16'h09CD
`define CUBE_LUT_2B32 16'h09D2
`define CUBE_LUT_2B34 16'h09D7
`define CUBE_LUT_2B37 16'h09DE
`define CUBE_LUT_2B39 16'h09E3
`define CUBE_LUT_2B3C 16'h09EA
`define CUBE_LUT_2B3E 16'h09EF
`define CUBE_LUT_2B41 16'h09F7
`define CUBE_LUT_2B43 16'h09FC
`define CUBE_LUT_2B46 16'h0A03
`define CUBE_LUT_2B48 16'h0A08
`define CUBE_LUT_2B4B 16'h0A10
`define CUBE_LUT_2B4D 16'h0A15
`define CUBE_LUT_2B4F 16'h0A1A
`define CUBE_LUT_2B52 16'h0A21
`define CUBE_LUT_2B54 16'h0A26
`define CUBE_LUT_2B57 16'h0A2E
`define CUBE_LUT_2B59 16'h0A33
`define CUBE_LUT_2B5C 16'h0A3A
`define CUBE_LUT_2B5E 16'h0A3F
`define CUBE_LUT_2B61 16'h0A47
`define CUBE_LUT_2B63 16'h0A4C
`define CUBE_LUT_2B66 16'h0A54
`define CUBE_LUT_2B68 16'h0A59
`define CUBE_LUT_2B6B 16'h0A61
`define CUBE_LUT_2B6D 16'h0A66
`define CUBE_LUT_2B6F 16'h0A6B
`define CUBE_LUT_2B72 16'h0A73
`define CUBE_LUT_2B74 16'h0A78
`define CUBE_LUT_2B77 16'h0A80
`define CUBE_LUT_2B79 16'h0A85
`define CUBE_LUT_2B7C 16'h0A8D
`define CUBE_LUT_2B7E 16'h0A92
`define CUBE_LUT_2B81 16'h0A9A
`define CUBE_LUT_2B83 16'h0A9F
`define CUBE_LUT_2B86 16'h0AA7
`define CUBE_LUT_2B88 16'h0AAD
`define CUBE_LUT_2B8A 16'h0AB2
`define CUBE_LUT_2B8D 16'h0ABA
`define CUBE_LUT_2B8F 16'h0ABF
`define CUBE_LUT_2B92 16'h0AC7
`define CUBE_LUT_2B94 16'h0ACD
`define CUBE_LUT_2B97 16'h0AD5
`define CUBE_LUT_2B99 16'h0ADA
`define CUBE_LUT_2B9C 16'h0AE2
`define CUBE_LUT_2B9E 16'h0AE8
`define CUBE_LUT_2BA1 16'h0AF0
`define CUBE_LUT_2BA3 16'h0AF5
`define CUBE_LUT_2BA6 16'h0AFE
`define CUBE_LUT_2BA8 16'h0B03
`define CUBE_LUT_2BAA 16'h0B09
`define CUBE_LUT_2BAD 16'h0B11
`define CUBE_LUT_2BAF 16'h0B16
`define CUBE_LUT_2BB2 16'h0B1F
`define CUBE_LUT_2BB4 16'h0B24
`define CUBE_LUT_2BB7 16'h0B2D
`define CUBE_LUT_2BB9 16'h0B32
`define CUBE_LUT_2BBC 16'h0B3B
`define CUBE_LUT_2BBE 16'h0B40
`define CUBE_LUT_2BC1 16'h0B49
`define CUBE_LUT_2BC3 16'h0B4E
`define CUBE_LUT_2BC5 16'h0B54
`define CUBE_LUT_2BC8 16'h0B5D
`define CUBE_LUT_2BCA 16'h0B62
`define CUBE_LUT_2BCD 16'h0B6B
`define CUBE_LUT_2BCF 16'h0B70
`define CUBE_LUT_2BD2 16'h0B79
`define CUBE_LUT_2BD4 16'h0B7F
`define CUBE_LUT_2BD7 16'h0B87
`define CUBE_LUT_2BD9 16'h0B8D
`define CUBE_LUT_2BDC 16'h0B96
`define CUBE_LUT_2BDE 16'h0B9C
`define CUBE_LUT_2BE0 16'h0BA1
`define CUBE_LUT_2BE3 16'h0BAA
`define CUBE_LUT_2BE5 16'h0BB0
`define CUBE_LUT_2BE8 16'h0BB9
`define CUBE_LUT_2BEA 16'h0BBF
`define CUBE_LUT_2BED 16'h0BC8
`define CUBE_LUT_2BEF 16'h0BCD
`define CUBE_LUT_2BF2 16'h0BD6
`define CUBE_LUT_2BF4 16'h0BDC
`define CUBE_LUT_2BF7 16'h0BE5
`define CUBE_LUT_2BF9 16'h0BEB
`define CUBE_LUT_2BFC 16'h0BF4
`define CUBE_LUT_2BFE 16'h0BFA
`define CUBE_LUT_2C00 16'h0C00
`define CUBE_LUT_2C01 16'h0C03
`define CUBE_LUT_2C03 16'h0C09
`define CUBE_LUT_2C04 16'h0C0C
`define CUBE_LUT_2C05 16'h0C0F
`define CUBE_LUT_2C06 16'h0C12
`define CUBE_LUT_2C08 16'h0C18
`define CUBE_LUT_2C09 16'h0C1B
`define CUBE_LUT_2C0A 16'h0C1E
`define CUBE_LUT_2C0B 16'h0C21
`define CUBE_LUT_2C0D 16'h0C27
`define CUBE_LUT_2C0E 16'h0C2B
`define CUBE_LUT_2C0F 16'h0C2E
`define CUBE_LUT_2C10 16'h0C31
`define CUBE_LUT_2C11 16'h0C34
`define CUBE_LUT_2C13 16'h0C3A
`define CUBE_LUT_2C14 16'h0C3D
`define CUBE_LUT_2C15 16'h0C40
`define CUBE_LUT_2C16 16'h0C43
`define CUBE_LUT_2C18 16'h0C4A
`define CUBE_LUT_2C19 16'h0C4D
`define CUBE_LUT_2C1A 16'h0C50
`define CUBE_LUT_2C1B 16'h0C53
`define CUBE_LUT_2C1C 16'h0C56
`define CUBE_LUT_2C1E 16'h0C5D
`define CUBE_LUT_2C1F 16'h0C60
`define CUBE_LUT_2C20 16'h0C63
`define CUBE_LUT_2C21 16'h0C66
`define CUBE_LUT_2C23 16'h0C6D
`define CUBE_LUT_2C24 16'h0C70
`define CUBE_LUT_2C25 16'h0C73
`define CUBE_LUT_2C26 16'h0C76
`define CUBE_LUT_2C28 16'h0C7D
`define CUBE_LUT_2C29 16'h0C80
`define CUBE_LUT_2C2A 16'h0C83
`define CUBE_LUT_2C2B 16'h0C86
`define CUBE_LUT_2C2C 16'h0C8A
`define CUBE_LUT_2C2E 16'h0C90
`define CUBE_LUT_2C2F 16'h0C94
`define CUBE_LUT_2C30 16'h0C97
`define CUBE_LUT_2C31 16'h0C9A
`define CUBE_LUT_2C33 16'h0CA1
`define CUBE_LUT_2C34 16'h0CA4
`define CUBE_LUT_2C35 16'h0CA7
`define CUBE_LUT_2C36 16'h0CAB
`define CUBE_LUT_2C38 16'h0CB1
`define CUBE_LUT_2C39 16'h0CB5
`define CUBE_LUT_2C3A 16'h0CB8
`define CUBE_LUT_2C3B 16'h0CBB
`define CUBE_LUT_2C3C 16'h0CBF
`define CUBE_LUT_2C3E 16'h0CC5
`define CUBE_LUT_2C3F 16'h0CC9
`define CUBE_LUT_2C40 16'h0CCC
`define CUBE_LUT_2C41 16'h0CD0
`define CUBE_LUT_2C43 16'h0CD6
`define CUBE_LUT_2C44 16'h0CDA
`define CUBE_LUT_2C45 16'h0CDD
`define CUBE_LUT_2C46 16'h0CE1
`define CUBE_LUT_2C47 16'h0CE4
`define CUBE_LUT_2C49 16'h0CEB
`define CUBE_LUT_2C4A 16'h0CEE
`define CUBE_LUT_2C4B 16'h0CF2
`define CUBE_LUT_2C4C 16'h0CF5
`define CUBE_LUT_2C4E 16'h0CFC
`define CUBE_LUT_2C4F 16'h0D00
`define CUBE_LUT_2C50 16'h0D03
`define CUBE_LUT_2C51 16'h0D07
`define CUBE_LUT_2C53 16'h0D0E
`define CUBE_LUT_2C54 16'h0D11
`define CUBE_LUT_2C55 16'h0D15
`define CUBE_LUT_2C56 16'h0D18
`define CUBE_LUT_2C57 16'h0D1C
`define CUBE_LUT_2C59 16'h0D23
`define CUBE_LUT_2C5A 16'h0D26
`define CUBE_LUT_2C5B 16'h0D2A
`define CUBE_LUT_2C5C 16'h0D2E
`define CUBE_LUT_2C5E 16'h0D35
`define CUBE_LUT_2C5F 16'h0D38
`define CUBE_LUT_2C60 16'h0D3C
`define CUBE_LUT_2C61 16'h0D3F
`define CUBE_LUT_2C63 16'h0D47
`define CUBE_LUT_2C64 16'h0D4A
`define CUBE_LUT_2C65 16'h0D4E
`define CUBE_LUT_2C66 16'h0D51
`define CUBE_LUT_2C67 16'h0D55
`define CUBE_LUT_2C69 16'h0D5C
`define CUBE_LUT_2C6A 16'h0D60
`define CUBE_LUT_2C6B 16'h0D64
`define CUBE_LUT_2C6C 16'h0D67
`define CUBE_LUT_2C6E 16'h0D6F
`define CUBE_LUT_2C6F 16'h0D72
`define CUBE_LUT_2C70 16'h0D76
`define CUBE_LUT_2C71 16'h0D7A
`define CUBE_LUT_2C72 16'h0D7D
`define CUBE_LUT_2C74 16'h0D85
`define CUBE_LUT_2C75 16'h0D89
`define CUBE_LUT_2C76 16'h0D8C
`define CUBE_LUT_2C77 16'h0D90
`define CUBE_LUT_2C79 16'h0D98
`define CUBE_LUT_2C7A 16'h0D9B
`define CUBE_LUT_2C7B 16'h0D9F
`define CUBE_LUT_2C7C 16'h0DA3
`define CUBE_LUT_2C7E 16'h0DAA
`define CUBE_LUT_2C7F 16'h0DAE
`define CUBE_LUT_2C80 16'h0DB2
`define CUBE_LUT_2C81 16'h0DB6
`define CUBE_LUT_2C82 16'h0DBA
`define CUBE_LUT_2C84 16'h0DC1
`define CUBE_LUT_2C85 16'h0DC5
`define CUBE_LUT_2C86 16'h0DC9
`define CUBE_LUT_2C87 16'h0DCD
`define CUBE_LUT_2C89 16'h0DD4
`define CUBE_LUT_2C8A 16'h0DD8
`define CUBE_LUT_2C8B 16'h0DDC
`define CUBE_LUT_2C8C 16'h0DE0
`define CUBE_LUT_2C8E 16'h0DE8
`define CUBE_LUT_2C8F 16'h0DEC
`define CUBE_LUT_2C90 16'h0DF0
`define CUBE_LUT_2C91 16'h0DF4
`define CUBE_LUT_2C92 16'h0DF7
`define CUBE_LUT_2C94 16'h0DFF
`define CUBE_LUT_2C95 16'h0E03
`define CUBE_LUT_2C96 16'h0E07
`define CUBE_LUT_2C97 16'h0E0B
`define CUBE_LUT_2C99 16'h0E13
`define CUBE_LUT_2C9A 16'h0E17
`define CUBE_LUT_2C9B 16'h0E1B
`define CUBE_LUT_2C9C 16'h0E1F
`define CUBE_LUT_2C9E 16'h0E27
`define CUBE_LUT_2C9F 16'h0E2B
`define CUBE_LUT_2CA0 16'h0E2F
`define CUBE_LUT_2CA1 16'h0E33
`define CUBE_LUT_2CA2 16'h0E37
`define CUBE_LUT_2CA4 16'h0E3F
`define CUBE_LUT_2CA5 16'h0E43
`define CUBE_LUT_2CA6 16'h0E47
`define CUBE_LUT_2CA7 16'h0E4B
`define CUBE_LUT_2CA9 16'h0E53
`define CUBE_LUT_2CAA 16'h0E57
`define CUBE_LUT_2CAB 16'h0E5B
`define CUBE_LUT_2CAC 16'h0E60
`define CUBE_LUT_2CAD 16'h0E64
`define CUBE_LUT_2CAF 16'h0E6C
`define CUBE_LUT_2CB0 16'h0E70
`define CUBE_LUT_2CB1 16'h0E74
`define CUBE_LUT_2CB2 16'h0E78
`define CUBE_LUT_2CB4 16'h0E80
`define CUBE_LUT_2CB5 16'h0E85
`define CUBE_LUT_2CB6 16'h0E89
`define CUBE_LUT_2CB7 16'h0E8D
`define CUBE_LUT_2CB9 16'h0E95
`define CUBE_LUT_2CBA 16'h0E99
`define CUBE_LUT_2CBB 16'h0E9E
`define CUBE_LUT_2CBC 16'h0EA2
`define CUBE_LUT_2CBD 16'h0EA6
`define CUBE_LUT_2CBF 16'h0EAF
`define CUBE_LUT_2CC0 16'h0EB3
`define CUBE_LUT_2CC1 16'h0EB7
`define CUBE_LUT_2CC2 16'h0EBB
`define CUBE_LUT_2CC4 16'h0EC4
`define CUBE_LUT_2CC5 16'h0EC8
`define CUBE_LUT_2CC6 16'h0ECC
`define CUBE_LUT_2CC7 16'h0ED1
`define CUBE_LUT_2CC9 16'h0ED9
`define CUBE_LUT_2CCA 16'h0EDD
`define CUBE_LUT_2CCB 16'h0EE2
`define CUBE_LUT_2CCC 16'h0EE6
`define CUBE_LUT_2CCD 16'h0EEA
`define CUBE_LUT_2CCF 16'h0EF3
`define CUBE_LUT_2CD0 16'h0EF7
`define CUBE_LUT_2CD1 16'h0EFC
`define CUBE_LUT_2CD2 16'h0F00
`define CUBE_LUT_2CD4 16'h0F09
`define CUBE_LUT_2CD5 16'h0F0D
`define CUBE_LUT_2CD6 16'h0F12
`define CUBE_LUT_2CD7 16'h0F16
`define CUBE_LUT_2CD8 16'h0F1A
`define CUBE_LUT_2CDA 16'h0F23
`define CUBE_LUT_2CDB 16'h0F28
`define CUBE_LUT_2CDC 16'h0F2C
`define CUBE_LUT_2CDD 16'h0F30
`define CUBE_LUT_2CDF 16'h0F39
`define CUBE_LUT_2CE0 16'h0F3E
`define CUBE_LUT_2CE1 16'h0F42
`define CUBE_LUT_2CE2 16'h0F47
`define CUBE_LUT_2CE4 16'h0F50
`define CUBE_LUT_2CE5 16'h0F54
`define CUBE_LUT_2CE6 16'h0F59
`define CUBE_LUT_2CE7 16'h0F5D
`define CUBE_LUT_2CE8 16'h0F62
`define CUBE_LUT_2CEA 16'h0F6B
`define CUBE_LUT_2CEB 16'h0F6F
`define CUBE_LUT_2CEC 16'h0F74
`define CUBE_LUT_2CED 16'h0F78
`define CUBE_LUT_2CEF 16'h0F81
`define CUBE_LUT_2CF0 16'h0F86
`define CUBE_LUT_2CF1 16'h0F8B
`define CUBE_LUT_2CF2 16'h0F8F
`define CUBE_LUT_2CF4 16'h0F98
`define CUBE_LUT_2CF5 16'h0F9D
`define CUBE_LUT_2CF6 16'h0FA1
`define CUBE_LUT_2CF7 16'h0FA6
`define CUBE_LUT_2CF8 16'h0FAB
`define CUBE_LUT_2CFA 16'h0FB4
`define CUBE_LUT_2CFB 16'h0FB9
`define CUBE_LUT_2CFC 16'h0FBD
`define CUBE_LUT_2CFD 16'h0FC2
`define CUBE_LUT_2CFF 16'h0FCB
`define CUBE_LUT_2D00 16'h0FD0
`define CUBE_LUT_2D01 16'h0FD5
`define CUBE_LUT_2D02 16'h0FD9
`define CUBE_LUT_2D03 16'h0FDE
`define CUBE_LUT_2D05 16'h0FE8
`define CUBE_LUT_2D06 16'h0FEC
`define CUBE_LUT_2D07 16'h0FF1
`define CUBE_LUT_2D08 16'h0FF6
`define CUBE_LUT_2D0A 16'h0FFF
`define CUBE_LUT_2D0B 16'h1002
`define CUBE_LUT_2D0C 16'h1004
`define CUBE_LUT_2D0D 16'h1007
`define CUBE_LUT_2D0F 16'h100C
`define CUBE_LUT_2D10 16'h100E
`define CUBE_LUT_2D11 16'h1010
`define CUBE_LUT_2D12 16'h1013
`define CUBE_LUT_2D13 16'h1015
`define CUBE_LUT_2D15 16'h101A
`define CUBE_LUT_2D16 16'h101C
`define CUBE_LUT_2D17 16'h101F
`define CUBE_LUT_2D18 16'h1021
`define CUBE_LUT_2D1A 16'h1026
`define CUBE_LUT_2D1B 16'h1029
`define CUBE_LUT_2D1C 16'h102B
`define CUBE_LUT_2D1D 16'h102E
`define CUBE_LUT_2D1F 16'h1032
`define CUBE_LUT_2D20 16'h1035
`define CUBE_LUT_2D21 16'h1037
`define CUBE_LUT_2D22 16'h103A
`define CUBE_LUT_2D23 16'h103C
`define CUBE_LUT_2D25 16'h1041
`define CUBE_LUT_2D26 16'h1044
`define CUBE_LUT_2D27 16'h1046
`define CUBE_LUT_2D28 16'h1049
`define CUBE_LUT_2D2A 16'h104E
`define CUBE_LUT_2D2B 16'h1050
`define CUBE_LUT_2D2C 16'h1053
`define CUBE_LUT_2D2D 16'h1055
`define CUBE_LUT_2D2F 16'h105A
`define CUBE_LUT_2D30 16'h105D
`define CUBE_LUT_2D31 16'h105F
`define CUBE_LUT_2D32 16'h1062
`define CUBE_LUT_2D33 16'h1064
`define CUBE_LUT_2D35 16'h1069
`define CUBE_LUT_2D36 16'h106C
`define CUBE_LUT_2D37 16'h106F
`define CUBE_LUT_2D38 16'h1071
`define CUBE_LUT_2D3A 16'h1076
`define CUBE_LUT_2D3B 16'h1079
`define CUBE_LUT_2D3C 16'h107B
`define CUBE_LUT_2D3D 16'h107E
`define CUBE_LUT_2D3E 16'h1080
`define CUBE_LUT_2D40 16'h1086
`define CUBE_LUT_2D41 16'h1088
`define CUBE_LUT_2D42 16'h108B
`define CUBE_LUT_2D43 16'h108D
`define CUBE_LUT_2D45 16'h1093
`define CUBE_LUT_2D46 16'h1095
`define CUBE_LUT_2D47 16'h1098
`define CUBE_LUT_2D48 16'h109A
`define CUBE_LUT_2D4A 16'h10A0
`define CUBE_LUT_2D4B 16'h10A2
`define CUBE_LUT_2D4C 16'h10A5
`define CUBE_LUT_2D4D 16'h10A8
`define CUBE_LUT_2D4E 16'h10AA
`define CUBE_LUT_2D50 16'h10AF
`define CUBE_LUT_2D51 16'h10B2
`define CUBE_LUT_2D52 16'h10B5
`define CUBE_LUT_2D53 16'h10B7
`define CUBE_LUT_2D55 16'h10BD
`define CUBE_LUT_2D56 16'h10BF
`define CUBE_LUT_2D57 16'h10C2
`define CUBE_LUT_2D58 16'h10C5
`define CUBE_LUT_2D5A 16'h10CA
`define CUBE_LUT_2D5B 16'h10CD
`define CUBE_LUT_2D5C 16'h10CF
`define CUBE_LUT_2D5D 16'h10D2
`define CUBE_LUT_2D5E 16'h10D5
`define CUBE_LUT_2D60 16'h10DA
`define CUBE_LUT_2D61 16'h10DD
`define CUBE_LUT_2D62 16'h10E0
`define CUBE_LUT_2D63 16'h10E2
`define CUBE_LUT_2D65 16'h10E8
`define CUBE_LUT_2D66 16'h10EB
`define CUBE_LUT_2D67 16'h10ED
`define CUBE_LUT_2D68 16'h10F0
`define CUBE_LUT_2D69 16'h10F3
`define CUBE_LUT_2D6B 16'h10F8
`define CUBE_LUT_2D6C 16'h10FB
`define CUBE_LUT_2D6D 16'h10FE
`define CUBE_LUT_2D6E 16'h1101
`define CUBE_LUT_2D70 16'h1106
`define CUBE_LUT_2D71 16'h1109
`define CUBE_LUT_2D72 16'h110C
`define CUBE_LUT_2D73 16'h110E
`define CUBE_LUT_2D75 16'h1114
`define CUBE_LUT_2D76 16'h1117
`define CUBE_LUT_2D77 16'h111A
`define CUBE_LUT_2D78 16'h111C
`define CUBE_LUT_2D79 16'h111F
`define CUBE_LUT_2D7B 16'h1125
`define CUBE_LUT_2D7C 16'h1128
`define CUBE_LUT_2D7D 16'h112B
`define CUBE_LUT_2D7E 16'h112D
`define CUBE_LUT_2D80 16'h1133
`define CUBE_LUT_2D81 16'h1136
`define CUBE_LUT_2D82 16'h1139
`define CUBE_LUT_2D83 16'h113C
`define CUBE_LUT_2D85 16'h1141
`define CUBE_LUT_2D86 16'h1144
`define CUBE_LUT_2D87 16'h1147
`define CUBE_LUT_2D88 16'h114A
`define CUBE_LUT_2D89 16'h114D
`define CUBE_LUT_2D8B 16'h1152
`define CUBE_LUT_2D8C 16'h1155
`define CUBE_LUT_2D8D 16'h1158
`define CUBE_LUT_2D8E 16'h115B
`define CUBE_LUT_2D90 16'h1161
`define CUBE_LUT_2D91 16'h1164
`define CUBE_LUT_2D92 16'h1167
`define CUBE_LUT_2D93 16'h116A
`define CUBE_LUT_2D94 16'h116D
`define CUBE_LUT_2D96 16'h1172
`define CUBE_LUT_2D97 16'h1175
`define CUBE_LUT_2D98 16'h1178
`define CUBE_LUT_2D99 16'h117B
`define CUBE_LUT_2D9B 16'h1181
`define CUBE_LUT_2D9C 16'h1184
`define CUBE_LUT_2D9D 16'h1187
`define CUBE_LUT_2D9E 16'h118A
`define CUBE_LUT_2DA0 16'h1190
`define CUBE_LUT_2DA1 16'h1193
`define CUBE_LUT_2DA2 16'h1196
`define CUBE_LUT_2DA3 16'h1199
`define CUBE_LUT_2DA4 16'h119C
`define CUBE_LUT_2DA6 16'h11A2
`define CUBE_LUT_2DA7 16'h11A5
`define CUBE_LUT_2DA8 16'h11A8
`define CUBE_LUT_2DA9 16'h11AB
`define CUBE_LUT_2DAB 16'h11B1
`define CUBE_LUT_2DAC 16'h11B4
`define CUBE_LUT_2DAD 16'h11B7
`define CUBE_LUT_2DAE 16'h11BA
`define CUBE_LUT_2DB0 16'h11C0
`define CUBE_LUT_2DB1 16'h11C3
`define CUBE_LUT_2DB2 16'h11C6
`define CUBE_LUT_2DB3 16'h11C9
`define CUBE_LUT_2DB4 16'h11CC
`define CUBE_LUT_2DB6 16'h11D2
`define CUBE_LUT_2DB7 16'h11D5
`define CUBE_LUT_2DB8 16'h11D8
`define CUBE_LUT_2DB9 16'h11DB
`define CUBE_LUT_2DBB 16'h11E1
`define CUBE_LUT_2DBC 16'h11E5
`define CUBE_LUT_2DBD 16'h11E8
`define CUBE_LUT_2DBE 16'h11EB
`define CUBE_LUT_2DC0 16'h11F1
`define CUBE_LUT_2DC1 16'h11F4
`define CUBE_LUT_2DC2 16'h11F7
`define CUBE_LUT_2DC3 16'h11FA
`define CUBE_LUT_2DC4 16'h11FD
`define CUBE_LUT_2DC6 16'h1204
`define CUBE_LUT_2DC7 16'h1207
`define CUBE_LUT_2DC8 16'h120A
`define CUBE_LUT_2DC9 16'h120D
`define CUBE_LUT_2DCB 16'h1213
`define CUBE_LUT_2DCC 16'h1216
`define CUBE_LUT_2DCD 16'h121A
`define CUBE_LUT_2DCE 16'h121D
`define CUBE_LUT_2DCF 16'h1220
`define CUBE_LUT_2DD1 16'h1226
`define CUBE_LUT_2DD2 16'h1229
`define CUBE_LUT_2DD3 16'h122D
`define CUBE_LUT_2DD4 16'h1230
`define CUBE_LUT_2DD6 16'h1236
`define CUBE_LUT_2DD7 16'h1239
`define CUBE_LUT_2DD8 16'h123C
`define CUBE_LUT_2DD9 16'h1240
`define CUBE_LUT_2DDB 16'h1246
`define CUBE_LUT_2DDC 16'h1249
`define CUBE_LUT_2DDD 16'h124D
`define CUBE_LUT_2DDE 16'h1250
`define CUBE_LUT_2DDF 16'h1253
`define CUBE_LUT_2DE1 16'h1259
`define CUBE_LUT_2DE2 16'h125D
`define CUBE_LUT_2DE3 16'h1260
`define CUBE_LUT_2DE4 16'h1263
`define CUBE_LUT_2DE6 16'h126A
`define CUBE_LUT_2DE7 16'h126D
`define CUBE_LUT_2DE8 16'h1270
`define CUBE_LUT_2DE9 16'h1274
`define CUBE_LUT_2DEB 16'h127A
`define CUBE_LUT_2DEC 16'h127D
`define CUBE_LUT_2DED 16'h1281
`define CUBE_LUT_2DEE 16'h1284
`define CUBE_LUT_2DEF 16'h1287
`define CUBE_LUT_2DF1 16'h128E
`define CUBE_LUT_2DF2 16'h1291
`define CUBE_LUT_2DF3 16'h1294
`define CUBE_LUT_2DF4 16'h1298
`define CUBE_LUT_2DF6 16'h129E
`define CUBE_LUT_2DF7 16'h12A2
`define CUBE_LUT_2DF8 16'h12A5
`define CUBE_LUT_2DF9 16'h12A8
`define CUBE_LUT_2DFA 16'h12AC
`define CUBE_LUT_2DFC 16'h12B3
`define CUBE_LUT_2DFD 16'h12B6
`define CUBE_LUT_2DFE 16'h12B9
`define CUBE_LUT_2DFF 16'h12BD
`define CUBE_LUT_2E01 16'h12C3
`define CUBE_LUT_2E02 16'h12C7
`define CUBE_LUT_2E03 16'h12CA
`define CUBE_LUT_2E04 16'h12CE
`define CUBE_LUT_2E06 16'h12D4
`define CUBE_LUT_2E07 16'h12D8
`define CUBE_LUT_2E08 16'h12DB
`define CUBE_LUT_2E09 16'h12DF
`define CUBE_LUT_2E0A 16'h12E2
`define CUBE_LUT_2E0C 16'h12E9
`define CUBE_LUT_2E0D 16'h12EC
`define CUBE_LUT_2E0E 16'h12F0
`define CUBE_LUT_2E0F 16'h12F3
`define CUBE_LUT_2E11 16'h12FA
`define CUBE_LUT_2E12 16'h12FD
`define CUBE_LUT_2E13 16'h1301
`define CUBE_LUT_2E14 16'h1304
`define CUBE_LUT_2E16 16'h130B
`define CUBE_LUT_2E17 16'h130F
`define CUBE_LUT_2E18 16'h1312
`define CUBE_LUT_2E19 16'h1316
`define CUBE_LUT_2E1A 16'h1319
`define CUBE_LUT_2E1C 16'h1320
`define CUBE_LUT_2E1D 16'h1324
`define CUBE_LUT_2E1E 16'h1327
`define CUBE_LUT_2E1F 16'h132B
`define CUBE_LUT_2E21 16'h1332
`define CUBE_LUT_2E22 16'h1335
`define CUBE_LUT_2E23 16'h1339
`define CUBE_LUT_2E24 16'h133C
`define CUBE_LUT_2E25 16'h1340
`define CUBE_LUT_2E27 16'h1347
`define CUBE_LUT_2E28 16'h134B
`define CUBE_LUT_2E29 16'h134E
`define CUBE_LUT_2E2A 16'h1352
`define CUBE_LUT_2E2C 16'h1359
`define CUBE_LUT_2E2D 16'h135C
`define CUBE_LUT_2E2E 16'h1360
`define CUBE_LUT_2E2F 16'h1364
`define CUBE_LUT_2E31 16'h136B
`define CUBE_LUT_2E32 16'h136E
`define CUBE_LUT_2E33 16'h1372
`define CUBE_LUT_2E34 16'h1376
`define CUBE_LUT_2E35 16'h1379
`define CUBE_LUT_2E37 16'h1380
`define CUBE_LUT_2E38 16'h1384
`define CUBE_LUT_2E39 16'h1388
`define CUBE_LUT_2E3A 16'h138B
`define CUBE_LUT_2E3C 16'h1393
`define CUBE_LUT_2E3D 16'h1396
`define CUBE_LUT_2E3E 16'h139A
`define CUBE_LUT_2E3F 16'h139D
`define CUBE_LUT_2E41 16'h13A5
`define CUBE_LUT_2E42 16'h13A8
`define CUBE_LUT_2E43 16'h13AC
`define CUBE_LUT_2E44 16'h13B0
`define CUBE_LUT_2E45 16'h13B3
`define CUBE_LUT_2E47 16'h13BB
`define CUBE_LUT_2E48 16'h13BF
`define CUBE_LUT_2E49 16'h13C2
`define CUBE_LUT_2E4A 16'h13C6
`define CUBE_LUT_2E4C 16'h13CD
`define CUBE_LUT_2E4D 16'h13D1
`define CUBE_LUT_2E4E 16'h13D5
`define CUBE_LUT_2E4F 16'h13D9
`define CUBE_LUT_2E51 16'h13E0
`define CUBE_LUT_2E52 16'h13E4
`define CUBE_LUT_2E53 16'h13E8
`define CUBE_LUT_2E54 16'h13EB
`define CUBE_LUT_2E55 16'h13EF
`define CUBE_LUT_2E57 16'h13F7
`define CUBE_LUT_2E58 16'h13FA
`define CUBE_LUT_2E59 16'h13FE
`define CUBE_LUT_2E5A 16'h1401
`define CUBE_LUT_2E5C 16'h1405
`define CUBE_LUT_2E5D 16'h1407
`define CUBE_LUT_2E5E 16'h1409
`define CUBE_LUT_2E5F 16'h140A
`define CUBE_LUT_2E60 16'h140C
`define CUBE_LUT_2E62 16'h1410
`define CUBE_LUT_2E63 16'h1412
`define CUBE_LUT_2E64 16'h1414
`define CUBE_LUT_2E65 16'h1416
`define CUBE_LUT_2E67 16'h141A
`define CUBE_LUT_2E68 16'h141C
`define CUBE_LUT_2E69 16'h141E
`define CUBE_LUT_2E6A 16'h1420
`define CUBE_LUT_2E6C 16'h1423
`define CUBE_LUT_2E6D 16'h1425
`define CUBE_LUT_2E6E 16'h1427
`define CUBE_LUT_2E6F 16'h1429
`define CUBE_LUT_2E70 16'h142B
`define CUBE_LUT_2E72 16'h142F
`define CUBE_LUT_2E73 16'h1431
`define CUBE_LUT_2E74 16'h1433
`define CUBE_LUT_2E75 16'h1435
`define CUBE_LUT_2E77 16'h1439
`define CUBE_LUT_2E78 16'h143B
`define CUBE_LUT_2E79 16'h143D
`define CUBE_LUT_2E7A 16'h143F
`define CUBE_LUT_2E7C 16'h1443
`define CUBE_LUT_2E7D 16'h1445
`define CUBE_LUT_2E7E 16'h1447
`define CUBE_LUT_2E7F 16'h1449
`define CUBE_LUT_2E80 16'h144A
`define CUBE_LUT_2E82 16'h144E
`define CUBE_LUT_2E83 16'h1450
`define CUBE_LUT_2E84 16'h1452
`define CUBE_LUT_2E85 16'h1454
`define CUBE_LUT_2E87 16'h1458
`define CUBE_LUT_2E88 16'h145A
`define CUBE_LUT_2E89 16'h145C
`define CUBE_LUT_2E8A 16'h145E
`define CUBE_LUT_2E8B 16'h1460
`define CUBE_LUT_2E8D 16'h1464
`define CUBE_LUT_2E8E 16'h1466
`define CUBE_LUT_2E8F 16'h1468
`define CUBE_LUT_2E90 16'h146A
`define CUBE_LUT_2E92 16'h146F
`define CUBE_LUT_2E93 16'h1471
`define CUBE_LUT_2E94 16'h1473
`define CUBE_LUT_2E95 16'h1475
`define CUBE_LUT_2E97 16'h1479
`define CUBE_LUT_2E98 16'h147B
`define CUBE_LUT_2E99 16'h147D
`define CUBE_LUT_2E9A 16'h147F
`define CUBE_LUT_2E9B 16'h1481
`define CUBE_LUT_2E9D 16'h1485
`define CUBE_LUT_2E9E 16'h1487
`define CUBE_LUT_2E9F 16'h1489
`define CUBE_LUT_2EA0 16'h148B
`define CUBE_LUT_2EA2 16'h148F
`define CUBE_LUT_2EA3 16'h1491
`define CUBE_LUT_2EA4 16'h1493
`define CUBE_LUT_2EA5 16'h1495
`define CUBE_LUT_2EA7 16'h149A
`define CUBE_LUT_2EA8 16'h149C
`define CUBE_LUT_2EA9 16'h149E
`define CUBE_LUT_2EAA 16'h14A0
`define CUBE_LUT_2EAB 16'h14A2
`define CUBE_LUT_2EAD 16'h14A6
`define CUBE_LUT_2EAE 16'h14A8
`define CUBE_LUT_2EAF 16'h14AA
`define CUBE_LUT_2EB0 16'h14AC
`define CUBE_LUT_2EB2 16'h14B1
`define CUBE_LUT_2EB3 16'h14B3
`define CUBE_LUT_2EB4 16'h14B5
`define CUBE_LUT_2EB5 16'h14B7
`define CUBE_LUT_2EB6 16'h14B9
`define CUBE_LUT_2EB8 16'h14BD
`define CUBE_LUT_2EB9 16'h14BF
`define CUBE_LUT_2EBA 16'h14C1
`define CUBE_LUT_2EBB 16'h14C4
`define CUBE_LUT_2EBD 16'h14C8
`define CUBE_LUT_2EBE 16'h14CA
`define CUBE_LUT_2EBF 16'h14CC
`define CUBE_LUT_2EC0 16'h14CE
`define CUBE_LUT_2EC2 16'h14D2
`define CUBE_LUT_2EC3 16'h14D5
`define CUBE_LUT_2EC4 16'h14D7
`define CUBE_LUT_2EC5 16'h14D9
`define CUBE_LUT_2EC6 16'h14DB
`define CUBE_LUT_2EC8 16'h14DF
`define CUBE_LUT_2EC9 16'h14E2
`define CUBE_LUT_2ECA 16'h14E4
`define CUBE_LUT_2ECB 16'h14E6
`define CUBE_LUT_2ECD 16'h14EA
`define CUBE_LUT_2ECE 16'h14EC
`define CUBE_LUT_2ECF 16'h14EF
`define CUBE_LUT_2ED0 16'h14F1
`define CUBE_LUT_2ED2 16'h14F5
`define CUBE_LUT_2ED3 16'h14F7
`define CUBE_LUT_2ED4 16'h14F9
`define CUBE_LUT_2ED5 16'h14FC
`define CUBE_LUT_2ED6 16'h14FE
`define CUBE_LUT_2ED8 16'h1502
`define CUBE_LUT_2ED9 16'h1504
`define CUBE_LUT_2EDA 16'h1507
`define CUBE_LUT_2EDB 16'h1509
`define CUBE_LUT_2EDD 16'h150D
`define CUBE_LUT_2EDE 16'h150F
`define CUBE_LUT_2EDF 16'h1512
`define CUBE_LUT_2EE0 16'h1514
`define CUBE_LUT_2EE2 16'h1518
`define CUBE_LUT_2EE3 16'h151A
`define CUBE_LUT_2EE4 16'h151D
`define CUBE_LUT_2EE5 16'h151F
`define CUBE_LUT_2EE6 16'h1521
`define CUBE_LUT_2EE8 16'h1526
`define CUBE_LUT_2EE9 16'h1528
`define CUBE_LUT_2EEA 16'h152A
`define CUBE_LUT_2EEB 16'h152C
`define CUBE_LUT_2EED 16'h1531
`define CUBE_LUT_2EEE 16'h1533
`define CUBE_LUT_2EEF 16'h1535
`define CUBE_LUT_2EF0 16'h1538
`define CUBE_LUT_2EF1 16'h153A
`define CUBE_LUT_2EF3 16'h153E
`define CUBE_LUT_2EF4 16'h1541
`define CUBE_LUT_2EF5 16'h1543
`define CUBE_LUT_2EF6 16'h1545
`define CUBE_LUT_2EF8 16'h154A
`define CUBE_LUT_2EF9 16'h154C
`define CUBE_LUT_2EFA 16'h154E
`define CUBE_LUT_2EFB 16'h1551
`define CUBE_LUT_2EFD 16'h1555
`define CUBE_LUT_2EFE 16'h1557
`define CUBE_LUT_2EFF 16'h155A
`define CUBE_LUT_2F00 16'h155C
`define CUBE_LUT_2F01 16'h155E
`define CUBE_LUT_2F03 16'h1563
`define CUBE_LUT_2F04 16'h1565
`define CUBE_LUT_2F05 16'h1568
`define CUBE_LUT_2F06 16'h156A
`define CUBE_LUT_2F08 16'h156E
`define CUBE_LUT_2F09 16'h1571
`define CUBE_LUT_2F0A 16'h1573
`define CUBE_LUT_2F0B 16'h1575
`define CUBE_LUT_2F0D 16'h157A
`define CUBE_LUT_2F0E 16'h157C
`define CUBE_LUT_2F0F 16'h157F
`define CUBE_LUT_2F10 16'h1581
`define CUBE_LUT_2F11 16'h1583
`define CUBE_LUT_2F13 16'h1588
`define CUBE_LUT_2F14 16'h158A
`define CUBE_LUT_2F15 16'h158D
`define CUBE_LUT_2F16 16'h158F
`define CUBE_LUT_2F18 16'h1594
`define CUBE_LUT_2F19 16'h1596
`define CUBE_LUT_2F1A 16'h1599
`define CUBE_LUT_2F1B 16'h159B
`define CUBE_LUT_2F1C 16'h159D
`define CUBE_LUT_2F1E 16'h15A2
`define CUBE_LUT_2F1F 16'h15A4
`define CUBE_LUT_2F20 16'h15A7
`define CUBE_LUT_2F21 16'h15A9
`define CUBE_LUT_2F23 16'h15AE
`define CUBE_LUT_2F24 16'h15B0
`define CUBE_LUT_2F25 16'h15B3
`define CUBE_LUT_2F26 16'h15B5
`define CUBE_LUT_2F28 16'h15BA
`define CUBE_LUT_2F29 16'h15BC
`define CUBE_LUT_2F2A 16'h15BF
`define CUBE_LUT_2F2B 16'h15C1
`define CUBE_LUT_2F2C 16'h15C4
`define CUBE_LUT_2F2E 16'h15C8
`define CUBE_LUT_2F2F 16'h15CB
`define CUBE_LUT_2F30 16'h15CD
`define CUBE_LUT_2F31 16'h15D0
`define CUBE_LUT_2F33 16'h15D5
`define CUBE_LUT_2F34 16'h15D7
`define CUBE_LUT_2F35 16'h15D9
`define CUBE_LUT_2F36 16'h15DC
`define CUBE_LUT_2F38 16'h15E1
`define CUBE_LUT_2F39 16'h15E3
`define CUBE_LUT_2F3A 16'h15E6
`define CUBE_LUT_2F3B 16'h15E8
`define CUBE_LUT_2F3C 16'h15EA
`define CUBE_LUT_2F3E 16'h15EF
`define CUBE_LUT_2F3F 16'h15F2
`define CUBE_LUT_2F40 16'h15F4
`define CUBE_LUT_2F41 16'h15F7
`define CUBE_LUT_2F43 16'h15FC
`define CUBE_LUT_2F44 16'h15FE
`define CUBE_LUT_2F45 16'h1601
`define CUBE_LUT_2F46 16'h1603
`define CUBE_LUT_2F47 16'h1606
`define CUBE_LUT_2F49 16'h160B
`define CUBE_LUT_2F4A 16'h160D
`define CUBE_LUT_2F4B 16'h1610
`define CUBE_LUT_2F4C 16'h1612
`define CUBE_LUT_2F4E 16'h1617
`define CUBE_LUT_2F4F 16'h161A
`define CUBE_LUT_2F50 16'h161C
`define CUBE_LUT_2F51 16'h161F
`define CUBE_LUT_2F53 16'h1624
`define CUBE_LUT_2F54 16'h1626
`define CUBE_LUT_2F55 16'h1629
`define CUBE_LUT_2F56 16'h162B
`define CUBE_LUT_2F57 16'h162E
`define CUBE_LUT_2F59 16'h1633
`define CUBE_LUT_2F5A 16'h1635
`define CUBE_LUT_2F5B 16'h1638
`define CUBE_LUT_2F5C 16'h163A
`define CUBE_LUT_2F5E 16'h163F
`define CUBE_LUT_2F5F 16'h1642
`define CUBE_LUT_2F60 16'h1645
`define CUBE_LUT_2F61 16'h1647
`define CUBE_LUT_2F63 16'h164C
`define CUBE_LUT_2F64 16'h164F
`define CUBE_LUT_2F65 16'h1651
`define CUBE_LUT_2F66 16'h1654
`define CUBE_LUT_2F67 16'h1656
`define CUBE_LUT_2F69 16'h165C
`define CUBE_LUT_2F6A 16'h165E
`define CUBE_LUT_2F6B 16'h1661
`define CUBE_LUT_2F6C 16'h1663
`define CUBE_LUT_2F6E 16'h1668
`define CUBE_LUT_2F6F 16'h166B
`define CUBE_LUT_2F70 16'h166E
`define CUBE_LUT_2F71 16'h1670
`define CUBE_LUT_2F73 16'h1675
`define CUBE_LUT_2F74 16'h1678
`define CUBE_LUT_2F75 16'h167B
`define CUBE_LUT_2F76 16'h167D
`define CUBE_LUT_2F77 16'h1680
`define CUBE_LUT_2F79 16'h1685
`define CUBE_LUT_2F7A 16'h1688
`define CUBE_LUT_2F7B 16'h168A
`define CUBE_LUT_2F7C 16'h168D
`define CUBE_LUT_2F7E 16'h1692
`define CUBE_LUT_2F7F 16'h1695
`define CUBE_LUT_2F80 16'h1698
`define CUBE_LUT_2F81 16'h169A
`define CUBE_LUT_2F82 16'h169D
`define CUBE_LUT_2F84 16'h16A2
`define CUBE_LUT_2F85 16'h16A5
`define CUBE_LUT_2F86 16'h16A7
`define CUBE_LUT_2F87 16'h16AA
`define CUBE_LUT_2F89 16'h16AF
`define CUBE_LUT_2F8A 16'h16B2
`define CUBE_LUT_2F8B 16'h16B5
`define CUBE_LUT_2F8C 16'h16B7
`define CUBE_LUT_2F8E 16'h16BD
`define CUBE_LUT_2F8F 16'h16BF
`define CUBE_LUT_2F90 16'h16C2
`define CUBE_LUT_2F91 16'h16C5
`define CUBE_LUT_2F92 16'h16C7
`define CUBE_LUT_2F94 16'h16CD
`define CUBE_LUT_2F95 16'h16CF
`define CUBE_LUT_2F96 16'h16D2
`define CUBE_LUT_2F97 16'h16D5
`define CUBE_LUT_2F99 16'h16DA
`define CUBE_LUT_2F9A 16'h16DD
`define CUBE_LUT_2F9B 16'h16E0
`define CUBE_LUT_2F9C 16'h16E2
`define CUBE_LUT_2F9E 16'h16E8
`define CUBE_LUT_2F9F 16'h16EB
`define CUBE_LUT_2FA0 16'h16ED
`define CUBE_LUT_2FA1 16'h16F0
`define CUBE_LUT_2FA2 16'h16F3
`define CUBE_LUT_2FA4 16'h16F8
`define CUBE_LUT_2FA5 16'h16FB
`define CUBE_LUT_2FA6 16'h16FE
`define CUBE_LUT_2FA7 16'h1700
`define CUBE_LUT_2FA9 16'h1706
`define CUBE_LUT_2FAA 16'h1709
`define CUBE_LUT_2FAB 16'h170B
`define CUBE_LUT_2FAC 16'h170E
`define CUBE_LUT_2FAD 16'h1711
`define CUBE_LUT_2FAF 16'h1716
`define CUBE_LUT_2FB0 16'h1719
`define CUBE_LUT_2FB1 16'h171C
`define CUBE_LUT_2FB2 16'h171F
`define CUBE_LUT_2FB4 16'h1724
`define CUBE_LUT_2FB5 16'h1727
`define CUBE_LUT_2FB6 16'h172A
`define CUBE_LUT_2FB7 16'h172D
`define CUBE_LUT_2FB9 16'h1732
`define CUBE_LUT_2FBA 16'h1735
`define CUBE_LUT_2FBB 16'h1738
`define CUBE_LUT_2FBC 16'h173B
`define CUBE_LUT_2FBD 16'h173E
`define CUBE_LUT_2FBF 16'h1743
`define CUBE_LUT_2FC0 16'h1746
`define CUBE_LUT_2FC1 16'h1749
`define CUBE_LUT_2FC2 16'h174C
`define CUBE_LUT_2FC4 16'h1751
`define CUBE_LUT_2FC5 16'h1754
`define CUBE_LUT_2FC6 16'h1757
`define CUBE_LUT_2FC7 16'h175A
`define CUBE_LUT_2FC9 16'h175F
`define CUBE_LUT_2FCA 16'h1762
`define CUBE_LUT_2FCB 16'h1765
`define CUBE_LUT_2FCC 16'h1768
`define CUBE_LUT_2FCD 16'h176B
`define CUBE_LUT_2FCF 16'h1770
`define CUBE_LUT_2FD0 16'h1773
`define CUBE_LUT_2FD1 16'h1776
`define CUBE_LUT_2FD2 16'h1779
`define CUBE_LUT_2FD4 16'h177F
`define CUBE_LUT_2FD5 16'h1782
`define CUBE_LUT_2FD6 16'h1785
`define CUBE_LUT_2FD7 16'h1787
`define CUBE_LUT_2FD8 16'h178A
`define CUBE_LUT_2FDA 16'h1790
`define CUBE_LUT_2FDB 16'h1793
`define CUBE_LUT_2FDC 16'h1796
`define CUBE_LUT_2FDD 16'h1799
`define CUBE_LUT_2FDF 16'h179F
`define CUBE_LUT_2FE0 16'h17A1
`define CUBE_LUT_2FE1 16'h17A4
`define CUBE_LUT_2FE2 16'h17A7
`define CUBE_LUT_2FE4 16'h17AD
`define CUBE_LUT_2FE5 16'h17B0
`define CUBE_LUT_2FE6 16'h17B3
`define CUBE_LUT_2FE7 16'h17B6
`define CUBE_LUT_2FE8 16'h17B9
`define CUBE_LUT_2FEA 16'h17BF
`define CUBE_LUT_2FEB 16'h17C2
`define CUBE_LUT_2FEC 16'h17C5
`define CUBE_LUT_2FED 16'h17C8
`define CUBE_LUT_2FEF 16'h17CD
`define CUBE_LUT_2FF0 16'h17D0
`define CUBE_LUT_2FF1 16'h17D3
`define CUBE_LUT_2FF2 16'h17D6
`define CUBE_LUT_2FF4 16'h17DC
`define CUBE_LUT_2FF5 16'h17DF
`define CUBE_LUT_2FF6 16'h17E2
`define CUBE_LUT_2FF7 16'h17E5
`define CUBE_LUT_2FF8 16'h17E8
`define CUBE_LUT_2FFA 16'h17EE
`define CUBE_LUT_2FFB 16'h17F1
`define CUBE_LUT_2FFC 16'h17F4
`define CUBE_LUT_2FFD 16'h17F7
`define CUBE_LUT_2FFF 16'h17FD
`define CUBE_LUT_3000 16'h1800
`define CUBE_LUT_3001 16'h1803
`define CUBE_LUT_3002 16'h1806
`define CUBE_LUT_3003 16'h1809
`define CUBE_LUT_3004 16'h180C
`define CUBE_LUT_3005 16'h180F
`define CUBE_LUT_3006 16'h1812
`define CUBE_LUT_3007 16'h1815
`define CUBE_LUT_3008 16'h1818
`define CUBE_LUT_3009 16'h181B
`define CUBE_LUT_300A 16'h181E
`define CUBE_LUT_300B 16'h1821
`define CUBE_LUT_300C 16'h1824
`define CUBE_LUT_300D 16'h1827
`define CUBE_LUT_300E 16'h182B
`define CUBE_LUT_300F 16'h182E
`define CUBE_LUT_3010 16'h1831
`define CUBE_LUT_3011 16'h1834
`define CUBE_LUT_3012 16'h1837
`define CUBE_LUT_3013 16'h183A
`define CUBE_LUT_3014 16'h183D
`define CUBE_LUT_3015 16'h1840
`define CUBE_LUT_3016 16'h1843
`define CUBE_LUT_3017 16'h1847
`define CUBE_LUT_3018 16'h184A
`define CUBE_LUT_3019 16'h184D
`define CUBE_LUT_301A 16'h1850
`define CUBE_LUT_301B 16'h1853
`define CUBE_LUT_301C 16'h1856
`define CUBE_LUT_301D 16'h1859
`define CUBE_LUT_301E 16'h185D
`define CUBE_LUT_301F 16'h1860
`define CUBE_LUT_3020 16'h1863
`define CUBE_LUT_3021 16'h1866
`define CUBE_LUT_3022 16'h1869
`define CUBE_LUT_3023 16'h186D
`define CUBE_LUT_3024 16'h1870
`define CUBE_LUT_3025 16'h1873
`define CUBE_LUT_3026 16'h1876
`define CUBE_LUT_3027 16'h187A
`define CUBE_LUT_3028 16'h187D
`define CUBE_LUT_3029 16'h1880
`define CUBE_LUT_302A 16'h1883
`define CUBE_LUT_302B 16'h1886
`define CUBE_LUT_302C 16'h188A
`define CUBE_LUT_302D 16'h188D
`define CUBE_LUT_302E 16'h1890
`define CUBE_LUT_302F 16'h1894
`define CUBE_LUT_3030 16'h1897
`define CUBE_LUT_3031 16'h189A
`define CUBE_LUT_3032 16'h189D
`define CUBE_LUT_3033 16'h18A1
`define CUBE_LUT_3034 16'h18A4
`define CUBE_LUT_3035 16'h18A7
`define CUBE_LUT_3036 16'h18AB
`define CUBE_LUT_3037 16'h18AE
`define CUBE_LUT_3038 16'h18B1
`define CUBE_LUT_3039 16'h18B5
`define CUBE_LUT_303A 16'h18B8
`define CUBE_LUT_303B 16'h18BB
`define CUBE_LUT_303C 16'h18BF
`define CUBE_LUT_303D 16'h18C2
`define CUBE_LUT_303E 16'h18C5
`define CUBE_LUT_303F 16'h18C9
`define CUBE_LUT_3040 16'h18CC
`define CUBE_LUT_3041 16'h18D0
`define CUBE_LUT_3042 16'h18D3
`define CUBE_LUT_3043 16'h18D6
`define CUBE_LUT_3044 16'h18DA
`define CUBE_LUT_3045 16'h18DD
`define CUBE_LUT_3046 16'h18E1
`define CUBE_LUT_3047 16'h18E4
`define CUBE_LUT_3048 16'h18E8
`define CUBE_LUT_3049 16'h18EB
`define CUBE_LUT_304A 16'h18EE
`define CUBE_LUT_304B 16'h18F2
`define CUBE_LUT_304C 16'h18F5
`define CUBE_LUT_304D 16'h18F9
`define CUBE_LUT_304E 16'h18FC
`define CUBE_LUT_304F 16'h1900
`define CUBE_LUT_3050 16'h1903
`define CUBE_LUT_3051 16'h1907
`define CUBE_LUT_3052 16'h190A
`define CUBE_LUT_3053 16'h190E
`define CUBE_LUT_3054 16'h1911
`define CUBE_LUT_3055 16'h1915
`define CUBE_LUT_3056 16'h1918
`define CUBE_LUT_3057 16'h191C
`define CUBE_LUT_3058 16'h191F
`define CUBE_LUT_3059 16'h1923
`define CUBE_LUT_305A 16'h1926
`define CUBE_LUT_305B 16'h192A
`define CUBE_LUT_305C 16'h192E
`define CUBE_LUT_305D 16'h1931
`define CUBE_LUT_305E 16'h1935
`define CUBE_LUT_305F 16'h1938
`define CUBE_LUT_3060 16'h193C
`define CUBE_LUT_3061 16'h193F
`define CUBE_LUT_3062 16'h1943
`define CUBE_LUT_3063 16'h1947
`define CUBE_LUT_3064 16'h194A
`define CUBE_LUT_3065 16'h194E
`define CUBE_LUT_3066 16'h1951
`define CUBE_LUT_3067 16'h1955
`define CUBE_LUT_3068 16'h1959
`define CUBE_LUT_3069 16'h195C
`define CUBE_LUT_306A 16'h1960
`define CUBE_LUT_306B 16'h1964
`define CUBE_LUT_306C 16'h1967
`define CUBE_LUT_306D 16'h196B
`define CUBE_LUT_306E 16'h196F
`define CUBE_LUT_306F 16'h1972
`define CUBE_LUT_3070 16'h1976
`define CUBE_LUT_3071 16'h197A
`define CUBE_LUT_3072 16'h197D
`define CUBE_LUT_3073 16'h1981
`define CUBE_LUT_3074 16'h1985
`define CUBE_LUT_3075 16'h1989
`define CUBE_LUT_3076 16'h198C
`define CUBE_LUT_3077 16'h1990
`define CUBE_LUT_3078 16'h1994
`define CUBE_LUT_3079 16'h1998
`define CUBE_LUT_307A 16'h199B
`define CUBE_LUT_307B 16'h199F
`define CUBE_LUT_307C 16'h19A3
`define CUBE_LUT_307D 16'h19A7
`define CUBE_LUT_307E 16'h19AA
`define CUBE_LUT_307F 16'h19AE
`define CUBE_LUT_3080 16'h19B2
`define CUBE_LUT_3081 16'h19B6
`define CUBE_LUT_3082 16'h19BA
`define CUBE_LUT_3083 16'h19BD
`define CUBE_LUT_3084 16'h19C1
`define CUBE_LUT_3085 16'h19C5
`define CUBE_LUT_3086 16'h19C9
`define CUBE_LUT_3087 16'h19CD
`define CUBE_LUT_3088 16'h19D1
`define CUBE_LUT_3089 16'h19D4
`define CUBE_LUT_308A 16'h19D8
`define CUBE_LUT_308B 16'h19DC
`define CUBE_LUT_308C 16'h19E0
`define CUBE_LUT_308D 16'h19E4
`define CUBE_LUT_308E 16'h19E8
`define CUBE_LUT_308F 16'h19EC
`define CUBE_LUT_3090 16'h19F0
`define CUBE_LUT_3091 16'h19F4
`define CUBE_LUT_3092 16'h19F7
`define CUBE_LUT_3093 16'h19FB
`define CUBE_LUT_3094 16'h19FF
`define CUBE_LUT_3095 16'h1A03
`define CUBE_LUT_3096 16'h1A07
`define CUBE_LUT_3097 16'h1A0B
`define CUBE_LUT_3098 16'h1A0F
`define CUBE_LUT_3099 16'h1A13
`define CUBE_LUT_309A 16'h1A17
`define CUBE_LUT_309B 16'h1A1B
`define CUBE_LUT_309C 16'h1A1F
`define CUBE_LUT_309D 16'h1A23
`define CUBE_LUT_309E 16'h1A27
`define CUBE_LUT_309F 16'h1A2B
`define CUBE_LUT_30A0 16'h1A2F
`define CUBE_LUT_30A1 16'h1A33
`define CUBE_LUT_30A2 16'h1A37
`define CUBE_LUT_30A3 16'h1A3B
`define CUBE_LUT_30A4 16'h1A3F
`define CUBE_LUT_30A5 16'h1A43
`define CUBE_LUT_30A6 16'h1A47
`define CUBE_LUT_30A7 16'h1A4B
`define CUBE_LUT_30A8 16'h1A4F
`define CUBE_LUT_30A9 16'h1A53
`define CUBE_LUT_30AA 16'h1A57
`define CUBE_LUT_30AB 16'h1A5B
`define CUBE_LUT_30AC 16'h1A60
`define CUBE_LUT_30AD 16'h1A64
`define CUBE_LUT_30AE 16'h1A68
`define CUBE_LUT_30AF 16'h1A6C
`define CUBE_LUT_30B0 16'h1A70
`define CUBE_LUT_30B1 16'h1A74
`define CUBE_LUT_30B2 16'h1A78
`define CUBE_LUT_30B3 16'h1A7C
`define CUBE_LUT_30B4 16'h1A80
`define CUBE_LUT_30B5 16'h1A85
`define CUBE_LUT_30B6 16'h1A89
`define CUBE_LUT_30B7 16'h1A8D
`define CUBE_LUT_30B8 16'h1A91
`define CUBE_LUT_30B9 16'h1A95
`define CUBE_LUT_30BA 16'h1A99
`define CUBE_LUT_30BB 16'h1A9E
`define CUBE_LUT_30BC 16'h1AA2
`define CUBE_LUT_30BD 16'h1AA6
`define CUBE_LUT_30BE 16'h1AAA
`define CUBE_LUT_30BF 16'h1AAF
`define CUBE_LUT_30C0 16'h1AB3
`define CUBE_LUT_30C1 16'h1AB7
`define CUBE_LUT_30C2 16'h1ABB
`define CUBE_LUT_30C3 16'h1ABF
`define CUBE_LUT_30C4 16'h1AC4
`define CUBE_LUT_30C5 16'h1AC8
`define CUBE_LUT_30C6 16'h1ACC
`define CUBE_LUT_30C7 16'h1AD1
`define CUBE_LUT_30C8 16'h1AD5
`define CUBE_LUT_30C9 16'h1AD9
`define CUBE_LUT_30CA 16'h1ADD
`define CUBE_LUT_30CB 16'h1AE2
`define CUBE_LUT_30CC 16'h1AE6
`define CUBE_LUT_30CD 16'h1AEA
`define CUBE_LUT_30CE 16'h1AEF
`define CUBE_LUT_30CF 16'h1AF3
`define CUBE_LUT_30D0 16'h1AF7
`define CUBE_LUT_30D1 16'h1AFC
`define CUBE_LUT_30D2 16'h1B00
`define CUBE_LUT_30D3 16'h1B04
`define CUBE_LUT_30D4 16'h1B09
`define CUBE_LUT_30D5 16'h1B0D
`define CUBE_LUT_30D6 16'h1B12
`define CUBE_LUT_30D7 16'h1B16
`define CUBE_LUT_30D8 16'h1B1A
`define CUBE_LUT_30D9 16'h1B1F
`define CUBE_LUT_30DA 16'h1B23
`define CUBE_LUT_30DB 16'h1B28
`define CUBE_LUT_30DC 16'h1B2C
`define CUBE_LUT_30DD 16'h1B30
`define CUBE_LUT_30DE 16'h1B35
`define CUBE_LUT_30DF 16'h1B39
`define CUBE_LUT_30E0 16'h1B3E
`define CUBE_LUT_30E1 16'h1B42
`define CUBE_LUT_30E2 16'h1B47
`define CUBE_LUT_30E3 16'h1B4B
`define CUBE_LUT_30E4 16'h1B50
`define CUBE_LUT_30E5 16'h1B54
`define CUBE_LUT_30E6 16'h1B59
`define CUBE_LUT_30E7 16'h1B5D
`define CUBE_LUT_30E8 16'h1B62
`define CUBE_LUT_30E9 16'h1B66
`define CUBE_LUT_30EA 16'h1B6B
`define CUBE_LUT_30EB 16'h1B6F
`define CUBE_LUT_30EC 16'h1B74
`define CUBE_LUT_30ED 16'h1B78
`define CUBE_LUT_30EE 16'h1B7D
`define CUBE_LUT_30EF 16'h1B81
`define CUBE_LUT_30F0 16'h1B86
`define CUBE_LUT_30F1 16'h1B8B
`define CUBE_LUT_30F2 16'h1B8F
`define CUBE_LUT_30F3 16'h1B94
`define CUBE_LUT_30F4 16'h1B98
`define CUBE_LUT_30F5 16'h1B9D
`define CUBE_LUT_30F6 16'h1BA1
`define CUBE_LUT_30F7 16'h1BA6
`define CUBE_LUT_30F8 16'h1BAB
`define CUBE_LUT_30F9 16'h1BAF
`define CUBE_LUT_30FA 16'h1BB4
`define CUBE_LUT_30FB 16'h1BB9
`define CUBE_LUT_30FC 16'h1BBD
`define CUBE_LUT_30FD 16'h1BC2
`define CUBE_LUT_30FE 16'h1BC7
`define CUBE_LUT_30FF 16'h1BCB
`define CUBE_LUT_3100 16'h1BD0
`define CUBE_LUT_3101 16'h1BD5
`define CUBE_LUT_3102 16'h1BD9
`define CUBE_LUT_3103 16'h1BDE
`define CUBE_LUT_3104 16'h1BE3
`define CUBE_LUT_3105 16'h1BE8
`define CUBE_LUT_3106 16'h1BEC
`define CUBE_LUT_3107 16'h1BF1
`define CUBE_LUT_3108 16'h1BF6
`define CUBE_LUT_3109 16'h1BFA
`define CUBE_LUT_310A 16'h1BFF
`define CUBE_LUT_310B 16'h1C02
`define CUBE_LUT_310C 16'h1C04
`define CUBE_LUT_310D 16'h1C07
`define CUBE_LUT_310E 16'h1C09
`define CUBE_LUT_310F 16'h1C0C
`define CUBE_LUT_3110 16'h1C0E
`define CUBE_LUT_3111 16'h1C10
`define CUBE_LUT_3112 16'h1C13
`define CUBE_LUT_3113 16'h1C15
`define CUBE_LUT_3114 16'h1C18
`define CUBE_LUT_3115 16'h1C1A
`define CUBE_LUT_3116 16'h1C1C
`define CUBE_LUT_3117 16'h1C1F
`define CUBE_LUT_3118 16'h1C21
`define CUBE_LUT_3119 16'h1C24
`define CUBE_LUT_311A 16'h1C26
`define CUBE_LUT_311B 16'h1C29
`define CUBE_LUT_311C 16'h1C2B
`define CUBE_LUT_311D 16'h1C2E
`define CUBE_LUT_311E 16'h1C30
`define CUBE_LUT_311F 16'h1C32
`define CUBE_LUT_3120 16'h1C35
`define CUBE_LUT_3121 16'h1C37
`define CUBE_LUT_3122 16'h1C3A
`define CUBE_LUT_3123 16'h1C3C
`define CUBE_LUT_3124 16'h1C3F
`define CUBE_LUT_3125 16'h1C41
`define CUBE_LUT_3126 16'h1C44
`define CUBE_LUT_3127 16'h1C46
`define CUBE_LUT_3128 16'h1C49
`define CUBE_LUT_3129 16'h1C4B
`define CUBE_LUT_312A 16'h1C4E
`define CUBE_LUT_312B 16'h1C50
`define CUBE_LUT_312C 16'h1C53
`define CUBE_LUT_312D 16'h1C55
`define CUBE_LUT_312E 16'h1C58
`define CUBE_LUT_312F 16'h1C5A
`define CUBE_LUT_3130 16'h1C5D
`define CUBE_LUT_3131 16'h1C5F
`define CUBE_LUT_3132 16'h1C62
`define CUBE_LUT_3133 16'h1C64
`define CUBE_LUT_3134 16'h1C67
`define CUBE_LUT_3135 16'h1C69
`define CUBE_LUT_3136 16'h1C6C
`define CUBE_LUT_3137 16'h1C6F
`define CUBE_LUT_3138 16'h1C71
`define CUBE_LUT_3139 16'h1C74
`define CUBE_LUT_313A 16'h1C76
`define CUBE_LUT_313B 16'h1C79
`define CUBE_LUT_313C 16'h1C7B
`define CUBE_LUT_313D 16'h1C7E
`define CUBE_LUT_313E 16'h1C80
`define CUBE_LUT_313F 16'h1C83
`define CUBE_LUT_3140 16'h1C86
`define CUBE_LUT_3141 16'h1C88
`define CUBE_LUT_3142 16'h1C8B
`define CUBE_LUT_3143 16'h1C8D
`define CUBE_LUT_3144 16'h1C90
`define CUBE_LUT_3145 16'h1C93
`define CUBE_LUT_3146 16'h1C95
`define CUBE_LUT_3147 16'h1C98
`define CUBE_LUT_3148 16'h1C9A
`define CUBE_LUT_3149 16'h1C9D
`define CUBE_LUT_314A 16'h1CA0
`define CUBE_LUT_314B 16'h1CA2
`define CUBE_LUT_314C 16'h1CA5
`define CUBE_LUT_314D 16'h1CA8
`define CUBE_LUT_314E 16'h1CAA
`define CUBE_LUT_314F 16'h1CAD
`define CUBE_LUT_3150 16'h1CAF
`define CUBE_LUT_3151 16'h1CB2
`define CUBE_LUT_3152 16'h1CB5
`define CUBE_LUT_3153 16'h1CB7
`define CUBE_LUT_3154 16'h1CBA
`define CUBE_LUT_3155 16'h1CBD
`define CUBE_LUT_3156 16'h1CBF
`define CUBE_LUT_3157 16'h1CC2
`define CUBE_LUT_3158 16'h1CC5
`define CUBE_LUT_3159 16'h1CC7
`define CUBE_LUT_315A 16'h1CCA
`define CUBE_LUT_315B 16'h1CCD
`define CUBE_LUT_315C 16'h1CCF
`define CUBE_LUT_315D 16'h1CD2
`define CUBE_LUT_315E 16'h1CD5
`define CUBE_LUT_315F 16'h1CD8
`define CUBE_LUT_3160 16'h1CDA
`define CUBE_LUT_3161 16'h1CDD
`define CUBE_LUT_3162 16'h1CE0
`define CUBE_LUT_3163 16'h1CE2
`define CUBE_LUT_3164 16'h1CE5
`define CUBE_LUT_3165 16'h1CE8
`define CUBE_LUT_3166 16'h1CEB
`define CUBE_LUT_3167 16'h1CED
`define CUBE_LUT_3168 16'h1CF0
`define CUBE_LUT_3169 16'h1CF3
`define CUBE_LUT_316A 16'h1CF6
`define CUBE_LUT_316B 16'h1CF8
`define CUBE_LUT_316C 16'h1CFB
`define CUBE_LUT_316D 16'h1CFE
`define CUBE_LUT_316E 16'h1D01
`define CUBE_LUT_316F 16'h1D03
`define CUBE_LUT_3170 16'h1D06
`define CUBE_LUT_3171 16'h1D09
`define CUBE_LUT_3172 16'h1D0C
`define CUBE_LUT_3173 16'h1D0E
`define CUBE_LUT_3174 16'h1D11
`define CUBE_LUT_3175 16'h1D14
`define CUBE_LUT_3176 16'h1D17
`define CUBE_LUT_3177 16'h1D1A
`define CUBE_LUT_3178 16'h1D1C
`define CUBE_LUT_3179 16'h1D1F
`define CUBE_LUT_317A 16'h1D22
`define CUBE_LUT_317B 16'h1D25
`define CUBE_LUT_317C 16'h1D28
`define CUBE_LUT_317D 16'h1D2B
`define CUBE_LUT_317E 16'h1D2D
`define CUBE_LUT_317F 16'h1D30
`define CUBE_LUT_3180 16'h1D33
`define CUBE_LUT_3181 16'h1D36
`define CUBE_LUT_3182 16'h1D39
`define CUBE_LUT_3183 16'h1D3C
`define CUBE_LUT_3184 16'h1D3E
`define CUBE_LUT_3185 16'h1D41
`define CUBE_LUT_3186 16'h1D44
`define CUBE_LUT_3187 16'h1D47
`define CUBE_LUT_3188 16'h1D4A
`define CUBE_LUT_3189 16'h1D4D
`define CUBE_LUT_318A 16'h1D50
`define CUBE_LUT_318B 16'h1D52
`define CUBE_LUT_318C 16'h1D55
`define CUBE_LUT_318D 16'h1D58
`define CUBE_LUT_318E 16'h1D5B
`define CUBE_LUT_318F 16'h1D5E
`define CUBE_LUT_3190 16'h1D61
`define CUBE_LUT_3191 16'h1D64
`define CUBE_LUT_3192 16'h1D67
`define CUBE_LUT_3193 16'h1D6A
`define CUBE_LUT_3194 16'h1D6D
`define CUBE_LUT_3195 16'h1D6F
`define CUBE_LUT_3196 16'h1D72
`define CUBE_LUT_3197 16'h1D75
`define CUBE_LUT_3198 16'h1D78
`define CUBE_LUT_3199 16'h1D7B
`define CUBE_LUT_319A 16'h1D7E
`define CUBE_LUT_319B 16'h1D81
`define CUBE_LUT_319C 16'h1D84
`define CUBE_LUT_319D 16'h1D87
`define CUBE_LUT_319E 16'h1D8A
`define CUBE_LUT_319F 16'h1D8D
`define CUBE_LUT_31A0 16'h1D90
`define CUBE_LUT_31A1 16'h1D93
`define CUBE_LUT_31A2 16'h1D96
`define CUBE_LUT_31A3 16'h1D99
`define CUBE_LUT_31A4 16'h1D9C
`define CUBE_LUT_31A5 16'h1D9F
`define CUBE_LUT_31A6 16'h1DA2
`define CUBE_LUT_31A7 16'h1DA5
`define CUBE_LUT_31A8 16'h1DA8
`define CUBE_LUT_31A9 16'h1DAB
`define CUBE_LUT_31AA 16'h1DAE
`define CUBE_LUT_31AB 16'h1DB1
`define CUBE_LUT_31AC 16'h1DB4
`define CUBE_LUT_31AD 16'h1DB7
`define CUBE_LUT_31AE 16'h1DBA
`define CUBE_LUT_31AF 16'h1DBD
`define CUBE_LUT_31B0 16'h1DC0
`define CUBE_LUT_31B1 16'h1DC3
`define CUBE_LUT_31B2 16'h1DC6
`define CUBE_LUT_31B3 16'h1DC9
`define CUBE_LUT_31B4 16'h1DCC
`define CUBE_LUT_31B5 16'h1DCF
`define CUBE_LUT_31B6 16'h1DD2
`define CUBE_LUT_31B7 16'h1DD5
`define CUBE_LUT_31B8 16'h1DD8
`define CUBE_LUT_31B9 16'h1DDB
`define CUBE_LUT_31BA 16'h1DDE
`define CUBE_LUT_31BB 16'h1DE1
`define CUBE_LUT_31BC 16'h1DE5
`define CUBE_LUT_31BD 16'h1DE8
`define CUBE_LUT_31BE 16'h1DEB
`define CUBE_LUT_31BF 16'h1DEE
`define CUBE_LUT_31C0 16'h1DF1
`define CUBE_LUT_31C1 16'h1DF4
`define CUBE_LUT_31C2 16'h1DF7
`define CUBE_LUT_31C3 16'h1DFA
`define CUBE_LUT_31C4 16'h1DFD
`define CUBE_LUT_31C5 16'h1E00
`define CUBE_LUT_31C6 16'h1E04
`define CUBE_LUT_31C7 16'h1E07
`define CUBE_LUT_31C8 16'h1E0A
`define CUBE_LUT_31C9 16'h1E0D
`define CUBE_LUT_31CA 16'h1E10
`define CUBE_LUT_31CB 16'h1E13
`define CUBE_LUT_31CC 16'h1E16
`define CUBE_LUT_31CD 16'h1E1A
`define CUBE_LUT_31CE 16'h1E1D
`define CUBE_LUT_31CF 16'h1E20
`define CUBE_LUT_31D0 16'h1E23
`define CUBE_LUT_31D1 16'h1E26
`define CUBE_LUT_31D2 16'h1E29
`define CUBE_LUT_31D3 16'h1E2D
`define CUBE_LUT_31D4 16'h1E30
`define CUBE_LUT_31D5 16'h1E33
`define CUBE_LUT_31D6 16'h1E36
`define CUBE_LUT_31D7 16'h1E39
`define CUBE_LUT_31D8 16'h1E3C
`define CUBE_LUT_31D9 16'h1E40
`define CUBE_LUT_31DA 16'h1E43
`define CUBE_LUT_31DB 16'h1E46
`define CUBE_LUT_31DC 16'h1E49
`define CUBE_LUT_31DD 16'h1E4D
`define CUBE_LUT_31DE 16'h1E50
`define CUBE_LUT_31DF 16'h1E53
`define CUBE_LUT_31E0 16'h1E56
`define CUBE_LUT_31E1 16'h1E59
`define CUBE_LUT_31E2 16'h1E5D
`define CUBE_LUT_31E3 16'h1E60
`define CUBE_LUT_31E4 16'h1E63
`define CUBE_LUT_31E5 16'h1E66
`define CUBE_LUT_31E6 16'h1E6A
`define CUBE_LUT_31E7 16'h1E6D
`define CUBE_LUT_31E8 16'h1E70
`define CUBE_LUT_31E9 16'h1E74
`define CUBE_LUT_31EA 16'h1E77
`define CUBE_LUT_31EB 16'h1E7A
`define CUBE_LUT_31EC 16'h1E7D
`define CUBE_LUT_31ED 16'h1E81
`define CUBE_LUT_31EE 16'h1E84
`define CUBE_LUT_31EF 16'h1E87
`define CUBE_LUT_31F0 16'h1E8B
`define CUBE_LUT_31F1 16'h1E8E
`define CUBE_LUT_31F2 16'h1E91
`define CUBE_LUT_31F3 16'h1E94
`define CUBE_LUT_31F4 16'h1E98
`define CUBE_LUT_31F5 16'h1E9B
`define CUBE_LUT_31F6 16'h1E9E
`define CUBE_LUT_31F7 16'h1EA2
`define CUBE_LUT_31F8 16'h1EA5
`define CUBE_LUT_31F9 16'h1EA8
`define CUBE_LUT_31FA 16'h1EAC
`define CUBE_LUT_31FB 16'h1EAF
`define CUBE_LUT_31FC 16'h1EB3
`define CUBE_LUT_31FD 16'h1EB6
`define CUBE_LUT_31FE 16'h1EB9
`define CUBE_LUT_31FF 16'h1EBD
`define CUBE_LUT_3200 16'h1EC0
`define CUBE_LUT_3201 16'h1EC3
`define CUBE_LUT_3202 16'h1EC7
`define CUBE_LUT_3203 16'h1ECA
`define CUBE_LUT_3204 16'h1ECE
`define CUBE_LUT_3205 16'h1ED1
`define CUBE_LUT_3206 16'h1ED4
`define CUBE_LUT_3207 16'h1ED8
`define CUBE_LUT_3208 16'h1EDB
`define CUBE_LUT_3209 16'h1EDF
`define CUBE_LUT_320A 16'h1EE2
`define CUBE_LUT_320B 16'h1EE5
`define CUBE_LUT_320C 16'h1EE9
`define CUBE_LUT_320D 16'h1EEC
`define CUBE_LUT_320E 16'h1EF0
`define CUBE_LUT_320F 16'h1EF3
`define CUBE_LUT_3210 16'h1EF7
`define CUBE_LUT_3211 16'h1EFA
`define CUBE_LUT_3212 16'h1EFD
`define CUBE_LUT_3213 16'h1F01
`define CUBE_LUT_3214 16'h1F04
`define CUBE_LUT_3215 16'h1F08
`define CUBE_LUT_3216 16'h1F0B
`define CUBE_LUT_3217 16'h1F0F
`define CUBE_LUT_3218 16'h1F12
`define CUBE_LUT_3219 16'h1F16
`define CUBE_LUT_321A 16'h1F19
`define CUBE_LUT_321B 16'h1F1D
`define CUBE_LUT_321C 16'h1F20
`define CUBE_LUT_321D 16'h1F24
`define CUBE_LUT_321E 16'h1F27
`define CUBE_LUT_321F 16'h1F2B
`define CUBE_LUT_3220 16'h1F2E
`define CUBE_LUT_3221 16'h1F32
`define CUBE_LUT_3222 16'h1F35
`define CUBE_LUT_3223 16'h1F39
`define CUBE_LUT_3224 16'h1F3C
`define CUBE_LUT_3225 16'h1F40
`define CUBE_LUT_3226 16'h1F43
`define CUBE_LUT_3227 16'h1F47
`define CUBE_LUT_3228 16'h1F4B
`define CUBE_LUT_3229 16'h1F4E
`define CUBE_LUT_322A 16'h1F52
`define CUBE_LUT_322B 16'h1F55
`define CUBE_LUT_322C 16'h1F59
`define CUBE_LUT_322D 16'h1F5C
`define CUBE_LUT_322E 16'h1F60
`define CUBE_LUT_322F 16'h1F64
`define CUBE_LUT_3230 16'h1F67
`define CUBE_LUT_3231 16'h1F6B
`define CUBE_LUT_3232 16'h1F6E
`define CUBE_LUT_3233 16'h1F72
`define CUBE_LUT_3234 16'h1F76
`define CUBE_LUT_3235 16'h1F79
`define CUBE_LUT_3236 16'h1F7D
`define CUBE_LUT_3237 16'h1F80
`define CUBE_LUT_3238 16'h1F84
`define CUBE_LUT_3239 16'h1F88
`define CUBE_LUT_323A 16'h1F8B
`define CUBE_LUT_323B 16'h1F8F
`define CUBE_LUT_323C 16'h1F93
`define CUBE_LUT_323D 16'h1F96
`define CUBE_LUT_323E 16'h1F9A
`define CUBE_LUT_323F 16'h1F9D
`define CUBE_LUT_3240 16'h1FA1
`define CUBE_LUT_3241 16'h1FA5
`define CUBE_LUT_3242 16'h1FA8
`define CUBE_LUT_3243 16'h1FAC
`define CUBE_LUT_3244 16'h1FB0
`define CUBE_LUT_3245 16'h1FB3
`define CUBE_LUT_3246 16'h1FB7
`define CUBE_LUT_3247 16'h1FBB
`define CUBE_LUT_3248 16'h1FBF
`define CUBE_LUT_3249 16'h1FC2
`define CUBE_LUT_324A 16'h1FC6
`define CUBE_LUT_324B 16'h1FCA
`define CUBE_LUT_324C 16'h1FCD
`define CUBE_LUT_324D 16'h1FD1
`define CUBE_LUT_324E 16'h1FD5
`define CUBE_LUT_324F 16'h1FD9
`define CUBE_LUT_3250 16'h1FDC
`define CUBE_LUT_3251 16'h1FE0
`define CUBE_LUT_3252 16'h1FE4
`define CUBE_LUT_3253 16'h1FE8
`define CUBE_LUT_3254 16'h1FEB
`define CUBE_LUT_3255 16'h1FEF
`define CUBE_LUT_3256 16'h1FF3
`define CUBE_LUT_3257 16'h1FF7
`define CUBE_LUT_3258 16'h1FFA
`define CUBE_LUT_3259 16'h1FFE
`define CUBE_LUT_325A 16'h2001
`define CUBE_LUT_325B 16'h2003
`define CUBE_LUT_325C 16'h2005
`define CUBE_LUT_325D 16'h2007
`define CUBE_LUT_325E 16'h2009
`define CUBE_LUT_325F 16'h200A
`define CUBE_LUT_3260 16'h200C
`define CUBE_LUT_3261 16'h200E
`define CUBE_LUT_3262 16'h2010
`define CUBE_LUT_3263 16'h2012
`define CUBE_LUT_3264 16'h2014
`define CUBE_LUT_3265 16'h2016
`define CUBE_LUT_3266 16'h2018
`define CUBE_LUT_3267 16'h201A
`define CUBE_LUT_3268 16'h201C
`define CUBE_LUT_3269 16'h201E
`define CUBE_LUT_326A 16'h2020
`define CUBE_LUT_326B 16'h2021
`define CUBE_LUT_326C 16'h2023
`define CUBE_LUT_326D 16'h2025
`define CUBE_LUT_326E 16'h2027
`define CUBE_LUT_326F 16'h2029
`define CUBE_LUT_3270 16'h202B
`define CUBE_LUT_3271 16'h202D
`define CUBE_LUT_3272 16'h202F
`define CUBE_LUT_3273 16'h2031
`define CUBE_LUT_3274 16'h2033
`define CUBE_LUT_3275 16'h2035
`define CUBE_LUT_3276 16'h2037
`define CUBE_LUT_3277 16'h2039
`define CUBE_LUT_3278 16'h203B
`define CUBE_LUT_3279 16'h203D
`define CUBE_LUT_327A 16'h203F
`define CUBE_LUT_327B 16'h2041
`define CUBE_LUT_327C 16'h2043
`define CUBE_LUT_327D 16'h2045
`define CUBE_LUT_327E 16'h2047
`define CUBE_LUT_327F 16'h2049
`define CUBE_LUT_3280 16'h204A
`define CUBE_LUT_3281 16'h204C
`define CUBE_LUT_3282 16'h204E
`define CUBE_LUT_3283 16'h2050
`define CUBE_LUT_3284 16'h2052
`define CUBE_LUT_3285 16'h2054
`define CUBE_LUT_3286 16'h2056
`define CUBE_LUT_3287 16'h2058
`define CUBE_LUT_3288 16'h205A
`define CUBE_LUT_3289 16'h205C
`define CUBE_LUT_328A 16'h205E
`define CUBE_LUT_328B 16'h2060
`define CUBE_LUT_328C 16'h2062
`define CUBE_LUT_328D 16'h2064
`define CUBE_LUT_328E 16'h2066
`define CUBE_LUT_328F 16'h2068
`define CUBE_LUT_3290 16'h206A
`define CUBE_LUT_3291 16'h206D
`define CUBE_LUT_3292 16'h206F
`define CUBE_LUT_3293 16'h2071
`define CUBE_LUT_3294 16'h2073
`define CUBE_LUT_3295 16'h2075
`define CUBE_LUT_3296 16'h2077
`define CUBE_LUT_3297 16'h2079
`define CUBE_LUT_3298 16'h207B
`define CUBE_LUT_3299 16'h207D
`define CUBE_LUT_329A 16'h207F
`define CUBE_LUT_329B 16'h2081
`define CUBE_LUT_329C 16'h2083
`define CUBE_LUT_329D 16'h2085
`define CUBE_LUT_329E 16'h2087
`define CUBE_LUT_329F 16'h2089
`define CUBE_LUT_32A0 16'h208B
`define CUBE_LUT_32A1 16'h208D
`define CUBE_LUT_32A2 16'h208F
`define CUBE_LUT_32A3 16'h2091
`define CUBE_LUT_32A4 16'h2093
`define CUBE_LUT_32A5 16'h2095
`define CUBE_LUT_32A6 16'h2097
`define CUBE_LUT_32A7 16'h209A
`define CUBE_LUT_32A8 16'h209C
`define CUBE_LUT_32A9 16'h209E
`define CUBE_LUT_32AA 16'h20A0
`define CUBE_LUT_32AB 16'h20A2
`define CUBE_LUT_32AC 16'h20A4
`define CUBE_LUT_32AD 16'h20A6
`define CUBE_LUT_32AE 16'h20A8
`define CUBE_LUT_32AF 16'h20AA
`define CUBE_LUT_32B0 16'h20AC
`define CUBE_LUT_32B1 16'h20AE
`define CUBE_LUT_32B2 16'h20B1
`define CUBE_LUT_32B3 16'h20B3
`define CUBE_LUT_32B4 16'h20B5
`define CUBE_LUT_32B5 16'h20B7
`define CUBE_LUT_32B6 16'h20B9
`define CUBE_LUT_32B7 16'h20BB
`define CUBE_LUT_32B8 16'h20BD
`define CUBE_LUT_32B9 16'h20BF
`define CUBE_LUT_32BA 16'h20C1
`define CUBE_LUT_32BB 16'h20C4
`define CUBE_LUT_32BC 16'h20C6
`define CUBE_LUT_32BD 16'h20C8
`define CUBE_LUT_32BE 16'h20CA
`define CUBE_LUT_32BF 16'h20CC
`define CUBE_LUT_32C0 16'h20CE
`define CUBE_LUT_32C1 16'h20D0
`define CUBE_LUT_32C2 16'h20D2
`define CUBE_LUT_32C3 16'h20D5
`define CUBE_LUT_32C4 16'h20D7
`define CUBE_LUT_32C5 16'h20D9
`define CUBE_LUT_32C6 16'h20DB
`define CUBE_LUT_32C7 16'h20DD
`define CUBE_LUT_32C8 16'h20DF
`define CUBE_LUT_32C9 16'h20E2
`define CUBE_LUT_32CA 16'h20E4
`define CUBE_LUT_32CB 16'h20E6
`define CUBE_LUT_32CC 16'h20E8
`define CUBE_LUT_32CD 16'h20EA
`define CUBE_LUT_32CE 16'h20EC
`define CUBE_LUT_32CF 16'h20EF
`define CUBE_LUT_32D0 16'h20F1
`define CUBE_LUT_32D1 16'h20F3
`define CUBE_LUT_32D2 16'h20F5
`define CUBE_LUT_32D3 16'h20F7
`define CUBE_LUT_32D4 16'h20F9
`define CUBE_LUT_32D5 16'h20FC
`define CUBE_LUT_32D6 16'h20FE
`define CUBE_LUT_32D7 16'h2100
`define CUBE_LUT_32D8 16'h2102
`define CUBE_LUT_32D9 16'h2104
`define CUBE_LUT_32DA 16'h2107
`define CUBE_LUT_32DB 16'h2109
`define CUBE_LUT_32DC 16'h210B
`define CUBE_LUT_32DD 16'h210D
`define CUBE_LUT_32DE 16'h210F
`define CUBE_LUT_32DF 16'h2112
`define CUBE_LUT_32E0 16'h2114
`define CUBE_LUT_32E1 16'h2116
`define CUBE_LUT_32E2 16'h2118
`define CUBE_LUT_32E3 16'h211A
`define CUBE_LUT_32E4 16'h211D
`define CUBE_LUT_32E5 16'h211F
`define CUBE_LUT_32E6 16'h2121
`define CUBE_LUT_32E7 16'h2123
`define CUBE_LUT_32E8 16'h2126
`define CUBE_LUT_32E9 16'h2128
`define CUBE_LUT_32EA 16'h212A
`define CUBE_LUT_32EB 16'h212C
`define CUBE_LUT_32EC 16'h212F
`define CUBE_LUT_32ED 16'h2131
`define CUBE_LUT_32EE 16'h2133
`define CUBE_LUT_32EF 16'h2135
`define CUBE_LUT_32F0 16'h2138
`define CUBE_LUT_32F1 16'h213A
`define CUBE_LUT_32F2 16'h213C
`define CUBE_LUT_32F3 16'h213E
`define CUBE_LUT_32F4 16'h2141
`define CUBE_LUT_32F5 16'h2143
`define CUBE_LUT_32F6 16'h2145
`define CUBE_LUT_32F7 16'h2147
`define CUBE_LUT_32F8 16'h214A
`define CUBE_LUT_32F9 16'h214C
`define CUBE_LUT_32FA 16'h214E
`define CUBE_LUT_32FB 16'h2151
`define CUBE_LUT_32FC 16'h2153
`define CUBE_LUT_32FD 16'h2155
`define CUBE_LUT_32FE 16'h2157
`define CUBE_LUT_32FF 16'h215A
`define CUBE_LUT_3300 16'h215C
`define CUBE_LUT_3301 16'h215E
`define CUBE_LUT_3302 16'h2161
`define CUBE_LUT_3303 16'h2163
`define CUBE_LUT_3304 16'h2165
`define CUBE_LUT_3305 16'h2168
`define CUBE_LUT_3306 16'h216A
`define CUBE_LUT_3307 16'h216C
`define CUBE_LUT_3308 16'h216E
`define CUBE_LUT_3309 16'h2171
`define CUBE_LUT_330A 16'h2173
`define CUBE_LUT_330B 16'h2175
`define CUBE_LUT_330C 16'h2178
`define CUBE_LUT_330D 16'h217A
`define CUBE_LUT_330E 16'h217C
`define CUBE_LUT_330F 16'h217F
`define CUBE_LUT_3310 16'h2181
`define CUBE_LUT_3311 16'h2183
`define CUBE_LUT_3312 16'h2186
`define CUBE_LUT_3313 16'h2188
`define CUBE_LUT_3314 16'h218A
`define CUBE_LUT_3315 16'h218D
`define CUBE_LUT_3316 16'h218F
`define CUBE_LUT_3317 16'h2192
`define CUBE_LUT_3318 16'h2194
`define CUBE_LUT_3319 16'h2196
`define CUBE_LUT_331A 16'h2199
`define CUBE_LUT_331B 16'h219B
`define CUBE_LUT_331C 16'h219D
`define CUBE_LUT_331D 16'h21A0
`define CUBE_LUT_331E 16'h21A2
`define CUBE_LUT_331F 16'h21A4
`define CUBE_LUT_3320 16'h21A7
`define CUBE_LUT_3321 16'h21A9
`define CUBE_LUT_3322 16'h21AC
`define CUBE_LUT_3323 16'h21AE
`define CUBE_LUT_3324 16'h21B0
`define CUBE_LUT_3325 16'h21B3
`define CUBE_LUT_3326 16'h21B5
`define CUBE_LUT_3327 16'h21B8
`define CUBE_LUT_3328 16'h21BA
`define CUBE_LUT_3329 16'h21BC
`define CUBE_LUT_332A 16'h21BF
`define CUBE_LUT_332B 16'h21C1
`define CUBE_LUT_332C 16'h21C4
`define CUBE_LUT_332D 16'h21C6
`define CUBE_LUT_332E 16'h21C8
`define CUBE_LUT_332F 16'h21CB
`define CUBE_LUT_3330 16'h21CD
`define CUBE_LUT_3331 16'h21D0
`define CUBE_LUT_3332 16'h21D2
`define CUBE_LUT_3333 16'h21D5
`define CUBE_LUT_3334 16'h21D7
`define CUBE_LUT_3335 16'h21D9
`define CUBE_LUT_3336 16'h21DC
`define CUBE_LUT_3337 16'h21DE
`define CUBE_LUT_3338 16'h21E1
`define CUBE_LUT_3339 16'h21E3
`define CUBE_LUT_333A 16'h21E6
`define CUBE_LUT_333B 16'h21E8
`define CUBE_LUT_333C 16'h21EA
`define CUBE_LUT_333D 16'h21ED
`define CUBE_LUT_333E 16'h21EF
`define CUBE_LUT_333F 16'h21F2
`define CUBE_LUT_3340 16'h21F4
`define CUBE_LUT_3341 16'h21F7
`define CUBE_LUT_3342 16'h21F9
`define CUBE_LUT_3343 16'h21FC
`define CUBE_LUT_3344 16'h21FE
`define CUBE_LUT_3345 16'h2201
`define CUBE_LUT_3346 16'h2203
`define CUBE_LUT_3347 16'h2206
`define CUBE_LUT_3348 16'h2208
`define CUBE_LUT_3349 16'h220B
`define CUBE_LUT_334A 16'h220D
`define CUBE_LUT_334B 16'h2210
`define CUBE_LUT_334C 16'h2212
`define CUBE_LUT_334D 16'h2215
`define CUBE_LUT_334E 16'h2217
`define CUBE_LUT_334F 16'h221A
`define CUBE_LUT_3350 16'h221C
`define CUBE_LUT_3351 16'h221F
`define CUBE_LUT_3352 16'h2221
`define CUBE_LUT_3353 16'h2224
`define CUBE_LUT_3354 16'h2226
`define CUBE_LUT_3355 16'h2229
`define CUBE_LUT_3356 16'h222B
`define CUBE_LUT_3357 16'h222E
`define CUBE_LUT_3358 16'h2230
`define CUBE_LUT_3359 16'h2233
`define CUBE_LUT_335A 16'h2235
`define CUBE_LUT_335B 16'h2238
`define CUBE_LUT_335C 16'h223A
`define CUBE_LUT_335D 16'h223D
`define CUBE_LUT_335E 16'h223F
`define CUBE_LUT_335F 16'h2242
`define CUBE_LUT_3360 16'h2245
`define CUBE_LUT_3361 16'h2247
`define CUBE_LUT_3362 16'h224A
`define CUBE_LUT_3363 16'h224C
`define CUBE_LUT_3364 16'h224F
`define CUBE_LUT_3365 16'h2251
`define CUBE_LUT_3366 16'h2254
`define CUBE_LUT_3367 16'h2256
`define CUBE_LUT_3368 16'h2259
`define CUBE_LUT_3369 16'h225C
`define CUBE_LUT_336A 16'h225E
`define CUBE_LUT_336B 16'h2261
`define CUBE_LUT_336C 16'h2263
`define CUBE_LUT_336D 16'h2266
`define CUBE_LUT_336E 16'h2268
`define CUBE_LUT_336F 16'h226B
`define CUBE_LUT_3370 16'h226E
`define CUBE_LUT_3371 16'h2270
`define CUBE_LUT_3372 16'h2273
`define CUBE_LUT_3373 16'h2275
`define CUBE_LUT_3374 16'h2278
`define CUBE_LUT_3375 16'h227B
`define CUBE_LUT_3376 16'h227D
`define CUBE_LUT_3377 16'h2280
`define CUBE_LUT_3378 16'h2282
`define CUBE_LUT_3379 16'h2285
`define CUBE_LUT_337A 16'h2288
`define CUBE_LUT_337B 16'h228A
`define CUBE_LUT_337C 16'h228D
`define CUBE_LUT_337D 16'h2290
`define CUBE_LUT_337E 16'h2292
`define CUBE_LUT_337F 16'h2295
`define CUBE_LUT_3380 16'h2298
`define CUBE_LUT_3381 16'h229A
`define CUBE_LUT_3382 16'h229D
`define CUBE_LUT_3383 16'h229F
`define CUBE_LUT_3384 16'h22A2
`define CUBE_LUT_3385 16'h22A5
`define CUBE_LUT_3386 16'h22A7
`define CUBE_LUT_3387 16'h22AA
`define CUBE_LUT_3388 16'h22AD
`define CUBE_LUT_3389 16'h22AF
`define CUBE_LUT_338A 16'h22B2
`define CUBE_LUT_338B 16'h22B5
`define CUBE_LUT_338C 16'h22B7
`define CUBE_LUT_338D 16'h22BA
`define CUBE_LUT_338E 16'h22BD
`define CUBE_LUT_338F 16'h22BF
`define CUBE_LUT_3390 16'h22C2
`define CUBE_LUT_3391 16'h22C5
`define CUBE_LUT_3392 16'h22C7
`define CUBE_LUT_3393 16'h22CA
`define CUBE_LUT_3394 16'h22CD
`define CUBE_LUT_3395 16'h22CF
`define CUBE_LUT_3396 16'h22D2
`define CUBE_LUT_3397 16'h22D5
`define CUBE_LUT_3398 16'h22D8
`define CUBE_LUT_3399 16'h22DA
`define CUBE_LUT_339A 16'h22DD
`define CUBE_LUT_339B 16'h22E0
`define CUBE_LUT_339C 16'h22E2
`define CUBE_LUT_339D 16'h22E5
`define CUBE_LUT_339E 16'h22E8
`define CUBE_LUT_339F 16'h22EB
`define CUBE_LUT_33A0 16'h22ED
`define CUBE_LUT_33A1 16'h22F0
`define CUBE_LUT_33A2 16'h22F3
`define CUBE_LUT_33A3 16'h22F5
`define CUBE_LUT_33A4 16'h22F8
`define CUBE_LUT_33A5 16'h22FB
`define CUBE_LUT_33A6 16'h22FE
`define CUBE_LUT_33A7 16'h2300
`define CUBE_LUT_33A8 16'h2303
`define CUBE_LUT_33A9 16'h2306
`define CUBE_LUT_33AA 16'h2309
`define CUBE_LUT_33AB 16'h230B
`define CUBE_LUT_33AC 16'h230E
`define CUBE_LUT_33AD 16'h2311
`define CUBE_LUT_33AE 16'h2314
`define CUBE_LUT_33AF 16'h2316
`define CUBE_LUT_33B0 16'h2319
`define CUBE_LUT_33B1 16'h231C
`define CUBE_LUT_33B2 16'h231F
`define CUBE_LUT_33B3 16'h2322
`define CUBE_LUT_33B4 16'h2324
`define CUBE_LUT_33B5 16'h2327
`define CUBE_LUT_33B6 16'h232A
`define CUBE_LUT_33B7 16'h232D
`define CUBE_LUT_33B8 16'h2330
`define CUBE_LUT_33B9 16'h2332
`define CUBE_LUT_33BA 16'h2335
`define CUBE_LUT_33BB 16'h2338
`define CUBE_LUT_33BC 16'h233B
`define CUBE_LUT_33BD 16'h233E
`define CUBE_LUT_33BE 16'h2340
`define CUBE_LUT_33BF 16'h2343
`define CUBE_LUT_33C0 16'h2346
`define CUBE_LUT_33C1 16'h2349
`define CUBE_LUT_33C2 16'h234C
`define CUBE_LUT_33C3 16'h234E
`define CUBE_LUT_33C4 16'h2351
`define CUBE_LUT_33C5 16'h2354
`define CUBE_LUT_33C6 16'h2357
`define CUBE_LUT_33C7 16'h235A
`define CUBE_LUT_33C8 16'h235D
`define CUBE_LUT_33C9 16'h235F
`define CUBE_LUT_33CA 16'h2362
`define CUBE_LUT_33CB 16'h2365
`define CUBE_LUT_33CC 16'h2368
`define CUBE_LUT_33CD 16'h236B
`define CUBE_LUT_33CE 16'h236E
`define CUBE_LUT_33CF 16'h2370
`define CUBE_LUT_33D0 16'h2373
`define CUBE_LUT_33D1 16'h2376
`define CUBE_LUT_33D2 16'h2379
`define CUBE_LUT_33D3 16'h237C
`define CUBE_LUT_33D4 16'h237F
`define CUBE_LUT_33D5 16'h2382
`define CUBE_LUT_33D6 16'h2385
`define CUBE_LUT_33D7 16'h2387
`define CUBE_LUT_33D8 16'h238A
`define CUBE_LUT_33D9 16'h238D
`define CUBE_LUT_33DA 16'h2390
`define CUBE_LUT_33DB 16'h2393
`define CUBE_LUT_33DC 16'h2396
`define CUBE_LUT_33DD 16'h2399
`define CUBE_LUT_33DE 16'h239C
`define CUBE_LUT_33DF 16'h239F
`define CUBE_LUT_33E0 16'h23A1
`define CUBE_LUT_33E1 16'h23A4
`define CUBE_LUT_33E2 16'h23A7
`define CUBE_LUT_33E3 16'h23AA
`define CUBE_LUT_33E4 16'h23AD
`define CUBE_LUT_33E5 16'h23B0
`define CUBE_LUT_33E6 16'h23B3
`define CUBE_LUT_33E7 16'h23B6
`define CUBE_LUT_33E8 16'h23B9
`define CUBE_LUT_33E9 16'h23BC
`define CUBE_LUT_33EA 16'h23BF
`define CUBE_LUT_33EB 16'h23C2
`define CUBE_LUT_33EC 16'h23C5
`define CUBE_LUT_33ED 16'h23C8
`define CUBE_LUT_33EE 16'h23CA
`define CUBE_LUT_33EF 16'h23CD
`define CUBE_LUT_33F0 16'h23D0
`define CUBE_LUT_33F1 16'h23D3
`define CUBE_LUT_33F2 16'h23D6
`define CUBE_LUT_33F3 16'h23D9
`define CUBE_LUT_33F4 16'h23DC
`define CUBE_LUT_33F5 16'h23DF
`define CUBE_LUT_33F6 16'h23E2
`define CUBE_LUT_33F7 16'h23E5
`define CUBE_LUT_33F8 16'h23E8
`define CUBE_LUT_33F9 16'h23EB
`define CUBE_LUT_33FA 16'h23EE
`define CUBE_LUT_33FB 16'h23F1
`define CUBE_LUT_33FC 16'h23F4
`define CUBE_LUT_33FD 16'h23F7
`define CUBE_LUT_33FE 16'h23FA
`define CUBE_LUT_33FF 16'h23FD
`define CUBE_LUT_3400 16'h2400
`define CUBE_LUT_3401 16'h2403
`define CUBE_LUT_3402 16'h2406
`define CUBE_LUT_3403 16'h2409
`define CUBE_LUT_3404 16'h240C
`define CUBE_LUT_3405 16'h240F
`define CUBE_LUT_3406 16'h2412
`define CUBE_LUT_3407 16'h2415
`define CUBE_LUT_3408 16'h2418
`define CUBE_LUT_3409 16'h241B
`define CUBE_LUT_340A 16'h241E
`define CUBE_LUT_340B 16'h2421
`define CUBE_LUT_340C 16'h2424
`define CUBE_LUT_340D 16'h2427
`define CUBE_LUT_340E 16'h242B
`define CUBE_LUT_340F 16'h242E
`define CUBE_LUT_3410 16'h2431
`define CUBE_LUT_3411 16'h2434
`define CUBE_LUT_3412 16'h2437
`define CUBE_LUT_3413 16'h243A
`define CUBE_LUT_3414 16'h243D
`define CUBE_LUT_3415 16'h2440
`define CUBE_LUT_3416 16'h2443
`define CUBE_LUT_3417 16'h2447
`define CUBE_LUT_3418 16'h244A
`define CUBE_LUT_3419 16'h244D
`define CUBE_LUT_341A 16'h2450
`define CUBE_LUT_341B 16'h2453
`define CUBE_LUT_341C 16'h2456
`define CUBE_LUT_341D 16'h2459
`define CUBE_LUT_341E 16'h245D
`define CUBE_LUT_341F 16'h2460
`define CUBE_LUT_3420 16'h2463
`define CUBE_LUT_3421 16'h2466
`define CUBE_LUT_3422 16'h2469
`define CUBE_LUT_3423 16'h246D
`define CUBE_LUT_3424 16'h2470
`define CUBE_LUT_3425 16'h2473
`define CUBE_LUT_3426 16'h2476
`define CUBE_LUT_3427 16'h247A
`define CUBE_LUT_3428 16'h247D
`define CUBE_LUT_3429 16'h2480
`define CUBE_LUT_342A 16'h2483
`define CUBE_LUT_342B 16'h2486
`define CUBE_LUT_342C 16'h248A
`define CUBE_LUT_342D 16'h248D
`define CUBE_LUT_342E 16'h2490
`define CUBE_LUT_342F 16'h2494
`define CUBE_LUT_3430 16'h2497
`define CUBE_LUT_3431 16'h249A
`define CUBE_LUT_3432 16'h249D
`define CUBE_LUT_3433 16'h24A1
`define CUBE_LUT_3434 16'h24A4
`define CUBE_LUT_3435 16'h24A7
`define CUBE_LUT_3436 16'h24AB
`define CUBE_LUT_3437 16'h24AE
`define CUBE_LUT_3438 16'h24B1
`define CUBE_LUT_3439 16'h24B5
`define CUBE_LUT_343A 16'h24B8
`define CUBE_LUT_343B 16'h24BB
`define CUBE_LUT_343C 16'h24BF
`define CUBE_LUT_343D 16'h24C2
`define CUBE_LUT_343E 16'h24C5
`define CUBE_LUT_343F 16'h24C9
`define CUBE_LUT_3440 16'h24CC
`define CUBE_LUT_3441 16'h24D0
`define CUBE_LUT_3442 16'h24D3
`define CUBE_LUT_3443 16'h24D6
`define CUBE_LUT_3444 16'h24DA
`define CUBE_LUT_3445 16'h24DD
`define CUBE_LUT_3446 16'h24E1
`define CUBE_LUT_3447 16'h24E4
`define CUBE_LUT_3448 16'h24E8
`define CUBE_LUT_3449 16'h24EB
`define CUBE_LUT_344A 16'h24EE
`define CUBE_LUT_344B 16'h24F2
`define CUBE_LUT_344C 16'h24F5
`define CUBE_LUT_344D 16'h24F9
`define CUBE_LUT_344E 16'h24FC
`define CUBE_LUT_344F 16'h2500
`define CUBE_LUT_3450 16'h2503
`define CUBE_LUT_3451 16'h2507
`define CUBE_LUT_3452 16'h250A
`define CUBE_LUT_3453 16'h250E
`define CUBE_LUT_3454 16'h2511
`define CUBE_LUT_3455 16'h2515
`define CUBE_LUT_3456 16'h2518
`define CUBE_LUT_3457 16'h251C
`define CUBE_LUT_3458 16'h251F
`define CUBE_LUT_3459 16'h2523
`define CUBE_LUT_345A 16'h2526
`define CUBE_LUT_345B 16'h252A
`define CUBE_LUT_345C 16'h252E
`define CUBE_LUT_345D 16'h2531
`define CUBE_LUT_345E 16'h2535
`define CUBE_LUT_345F 16'h2538
`define CUBE_LUT_3460 16'h253C
`define CUBE_LUT_3461 16'h253F
`define CUBE_LUT_3462 16'h2543
`define CUBE_LUT_3463 16'h2547
`define CUBE_LUT_3464 16'h254A
`define CUBE_LUT_3465 16'h254E
`define CUBE_LUT_3466 16'h2551
`define CUBE_LUT_3467 16'h2555
`define CUBE_LUT_3468 16'h2559
`define CUBE_LUT_3469 16'h255C
`define CUBE_LUT_346A 16'h2560
`define CUBE_LUT_346B 16'h2564
`define CUBE_LUT_346C 16'h2567
`define CUBE_LUT_346D 16'h256B
`define CUBE_LUT_346E 16'h256F
`define CUBE_LUT_346F 16'h2572
`define CUBE_LUT_3470 16'h2576
`define CUBE_LUT_3471 16'h257A
`define CUBE_LUT_3472 16'h257D
`define CUBE_LUT_3473 16'h2581
`define CUBE_LUT_3474 16'h2585
`define CUBE_LUT_3475 16'h2589
`define CUBE_LUT_3476 16'h258C
`define CUBE_LUT_3477 16'h2590
`define CUBE_LUT_3478 16'h2594
`define CUBE_LUT_3479 16'h2598
`define CUBE_LUT_347A 16'h259B
`define CUBE_LUT_347B 16'h259F
`define CUBE_LUT_347C 16'h25A3
`define CUBE_LUT_347D 16'h25A7
`define CUBE_LUT_347E 16'h25AA
`define CUBE_LUT_347F 16'h25AE
`define CUBE_LUT_3480 16'h25B2
`define CUBE_LUT_3481 16'h25B6
`define CUBE_LUT_3482 16'h25BA
`define CUBE_LUT_3483 16'h25BD
`define CUBE_LUT_3484 16'h25C1
`define CUBE_LUT_3485 16'h25C5
`define CUBE_LUT_3486 16'h25C9
`define CUBE_LUT_3487 16'h25CD
`define CUBE_LUT_3488 16'h25D1
`define CUBE_LUT_3489 16'h25D4
`define CUBE_LUT_348A 16'h25D8
`define CUBE_LUT_348B 16'h25DC
`define CUBE_LUT_348C 16'h25E0
`define CUBE_LUT_348D 16'h25E4
`define CUBE_LUT_348E 16'h25E8
`define CUBE_LUT_348F 16'h25EC
`define CUBE_LUT_3490 16'h25F0
`define CUBE_LUT_3491 16'h25F4
`define CUBE_LUT_3492 16'h25F7
`define CUBE_LUT_3493 16'h25FB
`define CUBE_LUT_3494 16'h25FF
`define CUBE_LUT_3495 16'h2603
`define CUBE_LUT_3496 16'h2607
`define CUBE_LUT_3497 16'h260B
`define CUBE_LUT_3498 16'h260F
`define CUBE_LUT_3499 16'h2613
`define CUBE_LUT_349A 16'h2617
`define CUBE_LUT_349B 16'h261B
`define CUBE_LUT_349C 16'h261F
`define CUBE_LUT_349D 16'h2623
`define CUBE_LUT_349E 16'h2627
`define CUBE_LUT_349F 16'h262B
`define CUBE_LUT_34A0 16'h262F
`define CUBE_LUT_34A1 16'h2633
`define CUBE_LUT_34A2 16'h2637
`define CUBE_LUT_34A3 16'h263B
`define CUBE_LUT_34A4 16'h263F
`define CUBE_LUT_34A5 16'h2643
`define CUBE_LUT_34A6 16'h2647
`define CUBE_LUT_34A7 16'h264B
`define CUBE_LUT_34A8 16'h264F
`define CUBE_LUT_34A9 16'h2653
`define CUBE_LUT_34AA 16'h2657
`define CUBE_LUT_34AB 16'h265B
`define CUBE_LUT_34AC 16'h2660
`define CUBE_LUT_34AD 16'h2664
`define CUBE_LUT_34AE 16'h2668
`define CUBE_LUT_34AF 16'h266C
`define CUBE_LUT_34B0 16'h2670
`define CUBE_LUT_34B1 16'h2674
`define CUBE_LUT_34B2 16'h2678
`define CUBE_LUT_34B3 16'h267C
`define CUBE_LUT_34B4 16'h2680
`define CUBE_LUT_34B5 16'h2685
`define CUBE_LUT_34B6 16'h2689
`define CUBE_LUT_34B7 16'h268D
`define CUBE_LUT_34B8 16'h2691
`define CUBE_LUT_34B9 16'h2695
`define CUBE_LUT_34BA 16'h2699
`define CUBE_LUT_34BB 16'h269E
`define CUBE_LUT_34BC 16'h26A2
`define CUBE_LUT_34BD 16'h26A6
`define CUBE_LUT_34BE 16'h26AA
`define CUBE_LUT_34BF 16'h26AF
`define CUBE_LUT_34C0 16'h26B3
`define CUBE_LUT_34C1 16'h26B7
`define CUBE_LUT_34C2 16'h26BB
`define CUBE_LUT_34C3 16'h26BF
`define CUBE_LUT_34C4 16'h26C4
`define CUBE_LUT_34C5 16'h26C8
`define CUBE_LUT_34C6 16'h26CC
`define CUBE_LUT_34C7 16'h26D1
`define CUBE_LUT_34C8 16'h26D5
`define CUBE_LUT_34C9 16'h26D9
`define CUBE_LUT_34CA 16'h26DD
`define CUBE_LUT_34CB 16'h26E2
`define CUBE_LUT_34CC 16'h26E6
`define CUBE_LUT_34CD 16'h26EA
`define CUBE_LUT_34CE 16'h26EF
`define CUBE_LUT_34CF 16'h26F3
`define CUBE_LUT_34D0 16'h26F7
`define CUBE_LUT_34D1 16'h26FC
`define CUBE_LUT_34D2 16'h2700
`define CUBE_LUT_34D3 16'h2704
`define CUBE_LUT_34D4 16'h2709
`define CUBE_LUT_34D5 16'h270D
`define CUBE_LUT_34D6 16'h2712
`define CUBE_LUT_34D7 16'h2716
`define CUBE_LUT_34D8 16'h271A
`define CUBE_LUT_34D9 16'h271F
`define CUBE_LUT_34DA 16'h2723
`define CUBE_LUT_34DB 16'h2728
`define CUBE_LUT_34DC 16'h272C
`define CUBE_LUT_34DD 16'h2730
`define CUBE_LUT_34DE 16'h2735
`define CUBE_LUT_34DF 16'h2739
`define CUBE_LUT_34E0 16'h273E
`define CUBE_LUT_34E1 16'h2742
`define CUBE_LUT_34E2 16'h2747
`define CUBE_LUT_34E3 16'h274B
`define CUBE_LUT_34E4 16'h2750
`define CUBE_LUT_34E5 16'h2754
`define CUBE_LUT_34E6 16'h2759
`define CUBE_LUT_34E7 16'h275D
`define CUBE_LUT_34E8 16'h2762
`define CUBE_LUT_34E9 16'h2766
`define CUBE_LUT_34EA 16'h276B
`define CUBE_LUT_34EB 16'h276F
`define CUBE_LUT_34EC 16'h2774
`define CUBE_LUT_34ED 16'h2778
`define CUBE_LUT_34EE 16'h277D
`define CUBE_LUT_34EF 16'h2781
`define CUBE_LUT_34F0 16'h2786
`define CUBE_LUT_34F1 16'h278B
`define CUBE_LUT_34F2 16'h278F
`define CUBE_LUT_34F3 16'h2794
`define CUBE_LUT_34F4 16'h2798
`define CUBE_LUT_34F5 16'h279D
`define CUBE_LUT_34F6 16'h27A1
`define CUBE_LUT_34F7 16'h27A6
`define CUBE_LUT_34F8 16'h27AB
`define CUBE_LUT_34F9 16'h27AF
`define CUBE_LUT_34FA 16'h27B4
`define CUBE_LUT_34FB 16'h27B9
`define CUBE_LUT_34FC 16'h27BD
`define CUBE_LUT_34FD 16'h27C2
`define CUBE_LUT_34FE 16'h27C7
`define CUBE_LUT_34FF 16'h27CB
`define CUBE_LUT_3500 16'h27D0
`define CUBE_LUT_3501 16'h27D5
`define CUBE_LUT_3502 16'h27D9
`define CUBE_LUT_3503 16'h27DE
`define CUBE_LUT_3504 16'h27E3
`define CUBE_LUT_3505 16'h27E8
`define CUBE_LUT_3506 16'h27EC
`define CUBE_LUT_3507 16'h27F1
`define CUBE_LUT_3508 16'h27F6
`define CUBE_LUT_3509 16'h27FA
`define CUBE_LUT_350A 16'h27FF
`define CUBE_LUT_350B 16'h2802
`define CUBE_LUT_350C 16'h2804
`define CUBE_LUT_350D 16'h2807
`define CUBE_LUT_350E 16'h2809
`define CUBE_LUT_350F 16'h280C
`define CUBE_LUT_3510 16'h280E
`define CUBE_LUT_3511 16'h2810
`define CUBE_LUT_3512 16'h2813
`define CUBE_LUT_3513 16'h2815
`define CUBE_LUT_3514 16'h2818
`define CUBE_LUT_3515 16'h281A
`define CUBE_LUT_3516 16'h281C
`define CUBE_LUT_3517 16'h281F
`define CUBE_LUT_3518 16'h2821
`define CUBE_LUT_3519 16'h2824
`define CUBE_LUT_351A 16'h2826
`define CUBE_LUT_351B 16'h2829
`define CUBE_LUT_351C 16'h282B
`define CUBE_LUT_351D 16'h282E
`define CUBE_LUT_351E 16'h2830
`define CUBE_LUT_351F 16'h2832
`define CUBE_LUT_3520 16'h2835
`define CUBE_LUT_3521 16'h2837
`define CUBE_LUT_3522 16'h283A
`define CUBE_LUT_3523 16'h283C
`define CUBE_LUT_3524 16'h283F
`define CUBE_LUT_3525 16'h2841
`define CUBE_LUT_3526 16'h2844
`define CUBE_LUT_3527 16'h2846
`define CUBE_LUT_3528 16'h2849
`define CUBE_LUT_3529 16'h284B
`define CUBE_LUT_352A 16'h284E
`define CUBE_LUT_352B 16'h2850
`define CUBE_LUT_352C 16'h2853
`define CUBE_LUT_352D 16'h2855
`define CUBE_LUT_352E 16'h2858
`define CUBE_LUT_352F 16'h285A
`define CUBE_LUT_3530 16'h285D
`define CUBE_LUT_3531 16'h285F
`define CUBE_LUT_3532 16'h2862
`define CUBE_LUT_3533 16'h2864
`define CUBE_LUT_3534 16'h2867
`define CUBE_LUT_3535 16'h2869
`define CUBE_LUT_3536 16'h286C
`define CUBE_LUT_3537 16'h286F
`define CUBE_LUT_3538 16'h2871
`define CUBE_LUT_3539 16'h2874
`define CUBE_LUT_353A 16'h2876
`define CUBE_LUT_353B 16'h2879
`define CUBE_LUT_353C 16'h287B
`define CUBE_LUT_353D 16'h287E
`define CUBE_LUT_353E 16'h2880
`define CUBE_LUT_353F 16'h2883
`define CUBE_LUT_3540 16'h2886
`define CUBE_LUT_3541 16'h2888
`define CUBE_LUT_3542 16'h288B
`define CUBE_LUT_3543 16'h288D
`define CUBE_LUT_3544 16'h2890
`define CUBE_LUT_3545 16'h2893
`define CUBE_LUT_3546 16'h2895
`define CUBE_LUT_3547 16'h2898
`define CUBE_LUT_3548 16'h289A
`define CUBE_LUT_3549 16'h289D
`define CUBE_LUT_354A 16'h28A0
`define CUBE_LUT_354B 16'h28A2
`define CUBE_LUT_354C 16'h28A5
`define CUBE_LUT_354D 16'h28A8
`define CUBE_LUT_354E 16'h28AA
`define CUBE_LUT_354F 16'h28AD
`define CUBE_LUT_3550 16'h28AF
`define CUBE_LUT_3551 16'h28B2
`define CUBE_LUT_3552 16'h28B5
`define CUBE_LUT_3553 16'h28B7
`define CUBE_LUT_3554 16'h28BA
`define CUBE_LUT_3555 16'h28BD
`define CUBE_LUT_3556 16'h28BF
`define CUBE_LUT_3557 16'h28C2
`define CUBE_LUT_3558 16'h28C5
`define CUBE_LUT_3559 16'h28C7
`define CUBE_LUT_355A 16'h28CA
`define CUBE_LUT_355B 16'h28CD
`define CUBE_LUT_355C 16'h28CF
`define CUBE_LUT_355D 16'h28D2
`define CUBE_LUT_355E 16'h28D5
`define CUBE_LUT_355F 16'h28D8
`define CUBE_LUT_3560 16'h28DA
`define CUBE_LUT_3561 16'h28DD
`define CUBE_LUT_3562 16'h28E0
`define CUBE_LUT_3563 16'h28E2
`define CUBE_LUT_3564 16'h28E5
`define CUBE_LUT_3565 16'h28E8
`define CUBE_LUT_3566 16'h28EB
`define CUBE_LUT_3567 16'h28ED
`define CUBE_LUT_3568 16'h28F0
`define CUBE_LUT_3569 16'h28F3
`define CUBE_LUT_356A 16'h28F6
`define CUBE_LUT_356B 16'h28F8
`define CUBE_LUT_356C 16'h28FB
`define CUBE_LUT_356D 16'h28FE
`define CUBE_LUT_356E 16'h2901
`define CUBE_LUT_356F 16'h2903
`define CUBE_LUT_3570 16'h2906
`define CUBE_LUT_3571 16'h2909
`define CUBE_LUT_3572 16'h290C
`define CUBE_LUT_3573 16'h290E
`define CUBE_LUT_3574 16'h2911
`define CUBE_LUT_3575 16'h2914
`define CUBE_LUT_3576 16'h2917
`define CUBE_LUT_3577 16'h291A
`define CUBE_LUT_3578 16'h291C
`define CUBE_LUT_3579 16'h291F
`define CUBE_LUT_357A 16'h2922
`define CUBE_LUT_357B 16'h2925
`define CUBE_LUT_357C 16'h2928
`define CUBE_LUT_357D 16'h292B
`define CUBE_LUT_357E 16'h292D
`define CUBE_LUT_357F 16'h2930
`define CUBE_LUT_3580 16'h2933
`define CUBE_LUT_3581 16'h2936
`define CUBE_LUT_3582 16'h2939
`define CUBE_LUT_3583 16'h293C
`define CUBE_LUT_3584 16'h293E
`define CUBE_LUT_3585 16'h2941
`define CUBE_LUT_3586 16'h2944
`define CUBE_LUT_3587 16'h2947
`define CUBE_LUT_3588 16'h294A
`define CUBE_LUT_3589 16'h294D
`define CUBE_LUT_358A 16'h2950
`define CUBE_LUT_358B 16'h2952
`define CUBE_LUT_358C 16'h2955
`define CUBE_LUT_358D 16'h2958
`define CUBE_LUT_358E 16'h295B
`define CUBE_LUT_358F 16'h295E
`define CUBE_LUT_3590 16'h2961
`define CUBE_LUT_3591 16'h2964
`define CUBE_LUT_3592 16'h2967
`define CUBE_LUT_3593 16'h296A
`define CUBE_LUT_3594 16'h296D
`define CUBE_LUT_3595 16'h296F
`define CUBE_LUT_3596 16'h2972
`define CUBE_LUT_3597 16'h2975
`define CUBE_LUT_3598 16'h2978
`define CUBE_LUT_3599 16'h297B
`define CUBE_LUT_359A 16'h297E
`define CUBE_LUT_359B 16'h2981
`define CUBE_LUT_359C 16'h2984
`define CUBE_LUT_359D 16'h2987
`define CUBE_LUT_359E 16'h298A
`define CUBE_LUT_359F 16'h298D
`define CUBE_LUT_35A0 16'h2990
`define CUBE_LUT_35A1 16'h2993
`define CUBE_LUT_35A2 16'h2996
`define CUBE_LUT_35A3 16'h2999
`define CUBE_LUT_35A4 16'h299C
`define CUBE_LUT_35A5 16'h299F
`define CUBE_LUT_35A6 16'h29A2
`define CUBE_LUT_35A7 16'h29A5
`define CUBE_LUT_35A8 16'h29A8
`define CUBE_LUT_35A9 16'h29AB
`define CUBE_LUT_35AA 16'h29AE
`define CUBE_LUT_35AB 16'h29B1
`define CUBE_LUT_35AC 16'h29B4
`define CUBE_LUT_35AD 16'h29B7
`define CUBE_LUT_35AE 16'h29BA
`define CUBE_LUT_35AF 16'h29BD
`define CUBE_LUT_35B0 16'h29C0
`define CUBE_LUT_35B1 16'h29C3
`define CUBE_LUT_35B2 16'h29C6
`define CUBE_LUT_35B3 16'h29C9
`define CUBE_LUT_35B4 16'h29CC
`define CUBE_LUT_35B5 16'h29CF
`define CUBE_LUT_35B6 16'h29D2
`define CUBE_LUT_35B7 16'h29D5
`define CUBE_LUT_35B8 16'h29D8
`define CUBE_LUT_35B9 16'h29DB
`define CUBE_LUT_35BA 16'h29DE
`define CUBE_LUT_35BB 16'h29E1
`define CUBE_LUT_35BC 16'h29E5
`define CUBE_LUT_35BD 16'h29E8
`define CUBE_LUT_35BE 16'h29EB
`define CUBE_LUT_35BF 16'h29EE
`define CUBE_LUT_35C0 16'h29F1
`define CUBE_LUT_35C1 16'h29F4
`define CUBE_LUT_35C2 16'h29F7
`define CUBE_LUT_35C3 16'h29FA
`define CUBE_LUT_35C4 16'h29FD
`define CUBE_LUT_35C5 16'h2A00
`define CUBE_LUT_35C6 16'h2A04
`define CUBE_LUT_35C7 16'h2A07
`define CUBE_LUT_35C8 16'h2A0A
`define CUBE_LUT_35C9 16'h2A0D
`define CUBE_LUT_35CA 16'h2A10
`define CUBE_LUT_35CB 16'h2A13
`define CUBE_LUT_35CC 16'h2A16
`define CUBE_LUT_35CD 16'h2A1A
`define CUBE_LUT_35CE 16'h2A1D
`define CUBE_LUT_35CF 16'h2A20
`define CUBE_LUT_35D0 16'h2A23
`define CUBE_LUT_35D1 16'h2A26
`define CUBE_LUT_35D2 16'h2A29
`define CUBE_LUT_35D3 16'h2A2D
`define CUBE_LUT_35D4 16'h2A30
`define CUBE_LUT_35D5 16'h2A33
`define CUBE_LUT_35D6 16'h2A36
`define CUBE_LUT_35D7 16'h2A39
`define CUBE_LUT_35D8 16'h2A3C
`define CUBE_LUT_35D9 16'h2A40
`define CUBE_LUT_35DA 16'h2A43
`define CUBE_LUT_35DB 16'h2A46
`define CUBE_LUT_35DC 16'h2A49
`define CUBE_LUT_35DD 16'h2A4D
`define CUBE_LUT_35DE 16'h2A50
`define CUBE_LUT_35DF 16'h2A53
`define CUBE_LUT_35E0 16'h2A56
`define CUBE_LUT_35E1 16'h2A59
`define CUBE_LUT_35E2 16'h2A5D
`define CUBE_LUT_35E3 16'h2A60
`define CUBE_LUT_35E4 16'h2A63
`define CUBE_LUT_35E5 16'h2A66
`define CUBE_LUT_35E6 16'h2A6A
`define CUBE_LUT_35E7 16'h2A6D
`define CUBE_LUT_35E8 16'h2A70
`define CUBE_LUT_35E9 16'h2A74
`define CUBE_LUT_35EA 16'h2A77
`define CUBE_LUT_35EB 16'h2A7A
`define CUBE_LUT_35EC 16'h2A7D
`define CUBE_LUT_35ED 16'h2A81
`define CUBE_LUT_35EE 16'h2A84
`define CUBE_LUT_35EF 16'h2A87
`define CUBE_LUT_35F0 16'h2A8B
`define CUBE_LUT_35F1 16'h2A8E
`define CUBE_LUT_35F2 16'h2A91
`define CUBE_LUT_35F3 16'h2A94
`define CUBE_LUT_35F4 16'h2A98
`define CUBE_LUT_35F5 16'h2A9B
`define CUBE_LUT_35F6 16'h2A9E
`define CUBE_LUT_35F7 16'h2AA2
`define CUBE_LUT_35F8 16'h2AA5
`define CUBE_LUT_35F9 16'h2AA8
`define CUBE_LUT_35FA 16'h2AAC
`define CUBE_LUT_35FB 16'h2AAF
`define CUBE_LUT_35FC 16'h2AB3
`define CUBE_LUT_35FD 16'h2AB6
`define CUBE_LUT_35FE 16'h2AB9
`define CUBE_LUT_35FF 16'h2ABD
`define CUBE_LUT_3600 16'h2AC0
`define CUBE_LUT_3601 16'h2AC3
`define CUBE_LUT_3602 16'h2AC7
`define CUBE_LUT_3603 16'h2ACA
`define CUBE_LUT_3604 16'h2ACE
`define CUBE_LUT_3605 16'h2AD1
`define CUBE_LUT_3606 16'h2AD4
`define CUBE_LUT_3607 16'h2AD8
`define CUBE_LUT_3608 16'h2ADB
`define CUBE_LUT_3609 16'h2ADF
`define CUBE_LUT_360A 16'h2AE2
`define CUBE_LUT_360B 16'h2AE5
`define CUBE_LUT_360C 16'h2AE9
`define CUBE_LUT_360D 16'h2AEC
`define CUBE_LUT_360E 16'h2AF0
`define CUBE_LUT_360F 16'h2AF3
`define CUBE_LUT_3610 16'h2AF7
`define CUBE_LUT_3611 16'h2AFA
`define CUBE_LUT_3612 16'h2AFD
`define CUBE_LUT_3613 16'h2B01
`define CUBE_LUT_3614 16'h2B04
`define CUBE_LUT_3615 16'h2B08
`define CUBE_LUT_3616 16'h2B0B
`define CUBE_LUT_3617 16'h2B0F
`define CUBE_LUT_3618 16'h2B12
`define CUBE_LUT_3619 16'h2B16
`define CUBE_LUT_361A 16'h2B19
`define CUBE_LUT_361B 16'h2B1D
`define CUBE_LUT_361C 16'h2B20
`define CUBE_LUT_361D 16'h2B24
`define CUBE_LUT_361E 16'h2B27
`define CUBE_LUT_361F 16'h2B2B
`define CUBE_LUT_3620 16'h2B2E
`define CUBE_LUT_3621 16'h2B32
`define CUBE_LUT_3622 16'h2B35
`define CUBE_LUT_3623 16'h2B39
`define CUBE_LUT_3624 16'h2B3C
`define CUBE_LUT_3625 16'h2B40
`define CUBE_LUT_3626 16'h2B43
`define CUBE_LUT_3627 16'h2B47
`define CUBE_LUT_3628 16'h2B4B
`define CUBE_LUT_3629 16'h2B4E
`define CUBE_LUT_362A 16'h2B52
`define CUBE_LUT_362B 16'h2B55
`define CUBE_LUT_362C 16'h2B59
`define CUBE_LUT_362D 16'h2B5C
`define CUBE_LUT_362E 16'h2B60
`define CUBE_LUT_362F 16'h2B64
`define CUBE_LUT_3630 16'h2B67
`define CUBE_LUT_3631 16'h2B6B
`define CUBE_LUT_3632 16'h2B6E
`define CUBE_LUT_3633 16'h2B72
`define CUBE_LUT_3634 16'h2B76
`define CUBE_LUT_3635 16'h2B79
`define CUBE_LUT_3636 16'h2B7D
`define CUBE_LUT_3637 16'h2B80
`define CUBE_LUT_3638 16'h2B84
`define CUBE_LUT_3639 16'h2B88
`define CUBE_LUT_363A 16'h2B8B
`define CUBE_LUT_363B 16'h2B8F
`define CUBE_LUT_363C 16'h2B93
`define CUBE_LUT_363D 16'h2B96
`define CUBE_LUT_363E 16'h2B9A
`define CUBE_LUT_363F 16'h2B9D
`define CUBE_LUT_3640 16'h2BA1
`define CUBE_LUT_3641 16'h2BA5
`define CUBE_LUT_3642 16'h2BA8
`define CUBE_LUT_3643 16'h2BAC
`define CUBE_LUT_3644 16'h2BB0
`define CUBE_LUT_3645 16'h2BB3
`define CUBE_LUT_3646 16'h2BB7
`define CUBE_LUT_3647 16'h2BBB
`define CUBE_LUT_3648 16'h2BBF
`define CUBE_LUT_3649 16'h2BC2
`define CUBE_LUT_364A 16'h2BC6
`define CUBE_LUT_364B 16'h2BCA
`define CUBE_LUT_364C 16'h2BCD
`define CUBE_LUT_364D 16'h2BD1
`define CUBE_LUT_364E 16'h2BD5
`define CUBE_LUT_364F 16'h2BD9
`define CUBE_LUT_3650 16'h2BDC
`define CUBE_LUT_3651 16'h2BE0
`define CUBE_LUT_3652 16'h2BE4
`define CUBE_LUT_3653 16'h2BE8
`define CUBE_LUT_3654 16'h2BEB
`define CUBE_LUT_3655 16'h2BEF
`define CUBE_LUT_3656 16'h2BF3
`define CUBE_LUT_3657 16'h2BF7
`define CUBE_LUT_3658 16'h2BFA
`define CUBE_LUT_3659 16'h2BFE
`define CUBE_LUT_365A 16'h2C01
`define CUBE_LUT_365B 16'h2C03
`define CUBE_LUT_365C 16'h2C05
`define CUBE_LUT_365D 16'h2C07
`define CUBE_LUT_365E 16'h2C09
`define CUBE_LUT_365F 16'h2C0A
`define CUBE_LUT_3660 16'h2C0C
`define CUBE_LUT_3661 16'h2C0E
`define CUBE_LUT_3662 16'h2C10
`define CUBE_LUT_3663 16'h2C12
`define CUBE_LUT_3664 16'h2C14
`define CUBE_LUT_3665 16'h2C16
`define CUBE_LUT_3666 16'h2C18
`define CUBE_LUT_3667 16'h2C1A
`define CUBE_LUT_3668 16'h2C1C
`define CUBE_LUT_3669 16'h2C1E
`define CUBE_LUT_366A 16'h2C20
`define CUBE_LUT_366B 16'h2C21
`define CUBE_LUT_366C 16'h2C23
`define CUBE_LUT_366D 16'h2C25
`define CUBE_LUT_366E 16'h2C27
`define CUBE_LUT_366F 16'h2C29
`define CUBE_LUT_3670 16'h2C2B
`define CUBE_LUT_3671 16'h2C2D
`define CUBE_LUT_3672 16'h2C2F
`define CUBE_LUT_3673 16'h2C31
`define CUBE_LUT_3674 16'h2C33
`define CUBE_LUT_3675 16'h2C35
`define CUBE_LUT_3676 16'h2C37
`define CUBE_LUT_3677 16'h2C39
`define CUBE_LUT_3678 16'h2C3B
`define CUBE_LUT_3679 16'h2C3D
`define CUBE_LUT_367A 16'h2C3F
`define CUBE_LUT_367B 16'h2C41
`define CUBE_LUT_367C 16'h2C43
`define CUBE_LUT_367D 16'h2C45
`define CUBE_LUT_367E 16'h2C47
`define CUBE_LUT_367F 16'h2C49
`define CUBE_LUT_3680 16'h2C4A
`define CUBE_LUT_3681 16'h2C4C
`define CUBE_LUT_3682 16'h2C4E
`define CUBE_LUT_3683 16'h2C50
`define CUBE_LUT_3684 16'h2C52
`define CUBE_LUT_3685 16'h2C54
`define CUBE_LUT_3686 16'h2C56
`define CUBE_LUT_3687 16'h2C58
`define CUBE_LUT_3688 16'h2C5A
`define CUBE_LUT_3689 16'h2C5C
`define CUBE_LUT_368A 16'h2C5E
`define CUBE_LUT_368B 16'h2C60
`define CUBE_LUT_368C 16'h2C62
`define CUBE_LUT_368D 16'h2C64
`define CUBE_LUT_368E 16'h2C66
`define CUBE_LUT_368F 16'h2C68
`define CUBE_LUT_3690 16'h2C6A
`define CUBE_LUT_3691 16'h2C6D
`define CUBE_LUT_3692 16'h2C6F
`define CUBE_LUT_3693 16'h2C71
`define CUBE_LUT_3694 16'h2C73
`define CUBE_LUT_3695 16'h2C75
`define CUBE_LUT_3696 16'h2C77
`define CUBE_LUT_3697 16'h2C79
`define CUBE_LUT_3698 16'h2C7B
`define CUBE_LUT_3699 16'h2C7D
`define CUBE_LUT_369A 16'h2C7F
`define CUBE_LUT_369B 16'h2C81
`define CUBE_LUT_369C 16'h2C83
`define CUBE_LUT_369D 16'h2C85
`define CUBE_LUT_369E 16'h2C87
`define CUBE_LUT_369F 16'h2C89
`define CUBE_LUT_36A0 16'h2C8B
`define CUBE_LUT_36A1 16'h2C8D
`define CUBE_LUT_36A2 16'h2C8F
`define CUBE_LUT_36A3 16'h2C91
`define CUBE_LUT_36A4 16'h2C93
`define CUBE_LUT_36A5 16'h2C95
`define CUBE_LUT_36A6 16'h2C97
`define CUBE_LUT_36A7 16'h2C9A
`define CUBE_LUT_36A8 16'h2C9C
`define CUBE_LUT_36A9 16'h2C9E
`define CUBE_LUT_36AA 16'h2CA0
`define CUBE_LUT_36AB 16'h2CA2
`define CUBE_LUT_36AC 16'h2CA4
`define CUBE_LUT_36AD 16'h2CA6
`define CUBE_LUT_36AE 16'h2CA8
`define CUBE_LUT_36AF 16'h2CAA
`define CUBE_LUT_36B0 16'h2CAC
`define CUBE_LUT_36B1 16'h2CAE
`define CUBE_LUT_36B2 16'h2CB1
`define CUBE_LUT_36B3 16'h2CB3
`define CUBE_LUT_36B4 16'h2CB5
`define CUBE_LUT_36B5 16'h2CB7
`define CUBE_LUT_36B6 16'h2CB9
`define CUBE_LUT_36B7 16'h2CBB
`define CUBE_LUT_36B8 16'h2CBD
`define CUBE_LUT_36B9 16'h2CBF
`define CUBE_LUT_36BA 16'h2CC1
`define CUBE_LUT_36BB 16'h2CC4
`define CUBE_LUT_36BC 16'h2CC6
`define CUBE_LUT_36BD 16'h2CC8
`define CUBE_LUT_36BE 16'h2CCA
`define CUBE_LUT_36BF 16'h2CCC
`define CUBE_LUT_36C0 16'h2CCE
`define CUBE_LUT_36C1 16'h2CD0
`define CUBE_LUT_36C2 16'h2CD2
`define CUBE_LUT_36C3 16'h2CD5
`define CUBE_LUT_36C4 16'h2CD7
`define CUBE_LUT_36C5 16'h2CD9
`define CUBE_LUT_36C6 16'h2CDB
`define CUBE_LUT_36C7 16'h2CDD
`define CUBE_LUT_36C8 16'h2CDF
`define CUBE_LUT_36C9 16'h2CE2
`define CUBE_LUT_36CA 16'h2CE4
`define CUBE_LUT_36CB 16'h2CE6
`define CUBE_LUT_36CC 16'h2CE8
`define CUBE_LUT_36CD 16'h2CEA
`define CUBE_LUT_36CE 16'h2CEC
`define CUBE_LUT_36CF 16'h2CEF
`define CUBE_LUT_36D0 16'h2CF1
`define CUBE_LUT_36D1 16'h2CF3
`define CUBE_LUT_36D2 16'h2CF5
`define CUBE_LUT_36D3 16'h2CF7
`define CUBE_LUT_36D4 16'h2CF9
`define CUBE_LUT_36D5 16'h2CFC
`define CUBE_LUT_36D6 16'h2CFE
`define CUBE_LUT_36D7 16'h2D00
`define CUBE_LUT_36D8 16'h2D02
`define CUBE_LUT_36D9 16'h2D04
`define CUBE_LUT_36DA 16'h2D07
`define CUBE_LUT_36DB 16'h2D09
`define CUBE_LUT_36DC 16'h2D0B
`define CUBE_LUT_36DD 16'h2D0D
`define CUBE_LUT_36DE 16'h2D0F
`define CUBE_LUT_36DF 16'h2D12
`define CUBE_LUT_36E0 16'h2D14
`define CUBE_LUT_36E1 16'h2D16
`define CUBE_LUT_36E2 16'h2D18
`define CUBE_LUT_36E3 16'h2D1A
`define CUBE_LUT_36E4 16'h2D1D
`define CUBE_LUT_36E5 16'h2D1F
`define CUBE_LUT_36E6 16'h2D21
`define CUBE_LUT_36E7 16'h2D23
`define CUBE_LUT_36E8 16'h2D26
`define CUBE_LUT_36E9 16'h2D28
`define CUBE_LUT_36EA 16'h2D2A
`define CUBE_LUT_36EB 16'h2D2C
`define CUBE_LUT_36EC 16'h2D2F
`define CUBE_LUT_36ED 16'h2D31
`define CUBE_LUT_36EE 16'h2D33
`define CUBE_LUT_36EF 16'h2D35
`define CUBE_LUT_36F0 16'h2D38
`define CUBE_LUT_36F1 16'h2D3A
`define CUBE_LUT_36F2 16'h2D3C
`define CUBE_LUT_36F3 16'h2D3E
`define CUBE_LUT_36F4 16'h2D41
`define CUBE_LUT_36F5 16'h2D43
`define CUBE_LUT_36F6 16'h2D45
`define CUBE_LUT_36F7 16'h2D47
`define CUBE_LUT_36F8 16'h2D4A
`define CUBE_LUT_36F9 16'h2D4C
`define CUBE_LUT_36FA 16'h2D4E
`define CUBE_LUT_36FB 16'h2D51
`define CUBE_LUT_36FC 16'h2D53
`define CUBE_LUT_36FD 16'h2D55
`define CUBE_LUT_36FE 16'h2D57
`define CUBE_LUT_36FF 16'h2D5A
`define CUBE_LUT_3700 16'h2D5C
`define CUBE_LUT_3701 16'h2D5E
`define CUBE_LUT_3702 16'h2D61
`define CUBE_LUT_3703 16'h2D63
`define CUBE_LUT_3704 16'h2D65
`define CUBE_LUT_3705 16'h2D68
`define CUBE_LUT_3706 16'h2D6A
`define CUBE_LUT_3707 16'h2D6C
`define CUBE_LUT_3708 16'h2D6E
`define CUBE_LUT_3709 16'h2D71
`define CUBE_LUT_370A 16'h2D73
`define CUBE_LUT_370B 16'h2D75
`define CUBE_LUT_370C 16'h2D78
`define CUBE_LUT_370D 16'h2D7A
`define CUBE_LUT_370E 16'h2D7C
`define CUBE_LUT_370F 16'h2D7F
`define CUBE_LUT_3710 16'h2D81
`define CUBE_LUT_3711 16'h2D83
`define CUBE_LUT_3712 16'h2D86
`define CUBE_LUT_3713 16'h2D88
`define CUBE_LUT_3714 16'h2D8A
`define CUBE_LUT_3715 16'h2D8D
`define CUBE_LUT_3716 16'h2D8F
`define CUBE_LUT_3717 16'h2D92
`define CUBE_LUT_3718 16'h2D94
`define CUBE_LUT_3719 16'h2D96
`define CUBE_LUT_371A 16'h2D99
`define CUBE_LUT_371B 16'h2D9B
`define CUBE_LUT_371C 16'h2D9D
`define CUBE_LUT_371D 16'h2DA0
`define CUBE_LUT_371E 16'h2DA2
`define CUBE_LUT_371F 16'h2DA4
`define CUBE_LUT_3720 16'h2DA7
`define CUBE_LUT_3721 16'h2DA9
`define CUBE_LUT_3722 16'h2DAC
`define CUBE_LUT_3723 16'h2DAE
`define CUBE_LUT_3724 16'h2DB0
`define CUBE_LUT_3725 16'h2DB3
`define CUBE_LUT_3726 16'h2DB5
`define CUBE_LUT_3727 16'h2DB8
`define CUBE_LUT_3728 16'h2DBA
`define CUBE_LUT_3729 16'h2DBC
`define CUBE_LUT_372A 16'h2DBF
`define CUBE_LUT_372B 16'h2DC1
`define CUBE_LUT_372C 16'h2DC4
`define CUBE_LUT_372D 16'h2DC6
`define CUBE_LUT_372E 16'h2DC8
`define CUBE_LUT_372F 16'h2DCB
`define CUBE_LUT_3730 16'h2DCD
`define CUBE_LUT_3731 16'h2DD0
`define CUBE_LUT_3732 16'h2DD2
`define CUBE_LUT_3733 16'h2DD5
`define CUBE_LUT_3734 16'h2DD7
`define CUBE_LUT_3735 16'h2DD9
`define CUBE_LUT_3736 16'h2DDC
`define CUBE_LUT_3737 16'h2DDE
`define CUBE_LUT_3738 16'h2DE1
`define CUBE_LUT_3739 16'h2DE3
`define CUBE_LUT_373A 16'h2DE6
`define CUBE_LUT_373B 16'h2DE8
`define CUBE_LUT_373C 16'h2DEA
`define CUBE_LUT_373D 16'h2DED
`define CUBE_LUT_373E 16'h2DEF
`define CUBE_LUT_373F 16'h2DF2
`define CUBE_LUT_3740 16'h2DF4
`define CUBE_LUT_3741 16'h2DF7
`define CUBE_LUT_3742 16'h2DF9
`define CUBE_LUT_3743 16'h2DFC
`define CUBE_LUT_3744 16'h2DFE
`define CUBE_LUT_3745 16'h2E01
`define CUBE_LUT_3746 16'h2E03
`define CUBE_LUT_3747 16'h2E06
`define CUBE_LUT_3748 16'h2E08
`define CUBE_LUT_3749 16'h2E0B
`define CUBE_LUT_374A 16'h2E0D
`define CUBE_LUT_374B 16'h2E10
`define CUBE_LUT_374C 16'h2E12
`define CUBE_LUT_374D 16'h2E15
`define CUBE_LUT_374E 16'h2E17
`define CUBE_LUT_374F 16'h2E1A
`define CUBE_LUT_3750 16'h2E1C
`define CUBE_LUT_3751 16'h2E1F
`define CUBE_LUT_3752 16'h2E21
`define CUBE_LUT_3753 16'h2E24
`define CUBE_LUT_3754 16'h2E26
`define CUBE_LUT_3755 16'h2E29
`define CUBE_LUT_3756 16'h2E2B
`define CUBE_LUT_3757 16'h2E2E
`define CUBE_LUT_3758 16'h2E30
`define CUBE_LUT_3759 16'h2E33
`define CUBE_LUT_375A 16'h2E35
`define CUBE_LUT_375B 16'h2E38
`define CUBE_LUT_375C 16'h2E3A
`define CUBE_LUT_375D 16'h2E3D
`define CUBE_LUT_375E 16'h2E3F
`define CUBE_LUT_375F 16'h2E42
`define CUBE_LUT_3760 16'h2E45
`define CUBE_LUT_3761 16'h2E47
`define CUBE_LUT_3762 16'h2E4A
`define CUBE_LUT_3763 16'h2E4C
`define CUBE_LUT_3764 16'h2E4F
`define CUBE_LUT_3765 16'h2E51
`define CUBE_LUT_3766 16'h2E54
`define CUBE_LUT_3767 16'h2E56
`define CUBE_LUT_3768 16'h2E59
`define CUBE_LUT_3769 16'h2E5C
`define CUBE_LUT_376A 16'h2E5E
`define CUBE_LUT_376B 16'h2E61
`define CUBE_LUT_376C 16'h2E63
`define CUBE_LUT_376D 16'h2E66
`define CUBE_LUT_376E 16'h2E68
`define CUBE_LUT_376F 16'h2E6B
`define CUBE_LUT_3770 16'h2E6E
`define CUBE_LUT_3771 16'h2E70
`define CUBE_LUT_3772 16'h2E73
`define CUBE_LUT_3773 16'h2E75
`define CUBE_LUT_3774 16'h2E78
`define CUBE_LUT_3775 16'h2E7B
`define CUBE_LUT_3776 16'h2E7D
`define CUBE_LUT_3777 16'h2E80
`define CUBE_LUT_3778 16'h2E82
`define CUBE_LUT_3779 16'h2E85
`define CUBE_LUT_377A 16'h2E88
`define CUBE_LUT_377B 16'h2E8A
`define CUBE_LUT_377C 16'h2E8D
`define CUBE_LUT_377D 16'h2E90
`define CUBE_LUT_377E 16'h2E92
`define CUBE_LUT_377F 16'h2E95
`define CUBE_LUT_3780 16'h2E98
`define CUBE_LUT_3781 16'h2E9A
`define CUBE_LUT_3782 16'h2E9D
`define CUBE_LUT_3783 16'h2E9F
`define CUBE_LUT_3784 16'h2EA2
`define CUBE_LUT_3785 16'h2EA5
`define CUBE_LUT_3786 16'h2EA7
`define CUBE_LUT_3787 16'h2EAA
`define CUBE_LUT_3788 16'h2EAD
`define CUBE_LUT_3789 16'h2EAF
`define CUBE_LUT_378A 16'h2EB2
`define CUBE_LUT_378B 16'h2EB5
`define CUBE_LUT_378C 16'h2EB7
`define CUBE_LUT_378D 16'h2EBA
`define CUBE_LUT_378E 16'h2EBD
`define CUBE_LUT_378F 16'h2EBF
`define CUBE_LUT_3790 16'h2EC2
`define CUBE_LUT_3791 16'h2EC5
`define CUBE_LUT_3792 16'h2EC7
`define CUBE_LUT_3793 16'h2ECA
`define CUBE_LUT_3794 16'h2ECD
`define CUBE_LUT_3795 16'h2ECF
`define CUBE_LUT_3796 16'h2ED2
`define CUBE_LUT_3797 16'h2ED5
`define CUBE_LUT_3798 16'h2ED8
`define CUBE_LUT_3799 16'h2EDA
`define CUBE_LUT_379A 16'h2EDD
`define CUBE_LUT_379B 16'h2EE0
`define CUBE_LUT_379C 16'h2EE2
`define CUBE_LUT_379D 16'h2EE5
`define CUBE_LUT_379E 16'h2EE8
`define CUBE_LUT_379F 16'h2EEB
`define CUBE_LUT_37A0 16'h2EED
`define CUBE_LUT_37A1 16'h2EF0
`define CUBE_LUT_37A2 16'h2EF3
`define CUBE_LUT_37A3 16'h2EF5
`define CUBE_LUT_37A4 16'h2EF8
`define CUBE_LUT_37A5 16'h2EFB
`define CUBE_LUT_37A6 16'h2EFE
`define CUBE_LUT_37A7 16'h2F00
`define CUBE_LUT_37A8 16'h2F03
`define CUBE_LUT_37A9 16'h2F06
`define CUBE_LUT_37AA 16'h2F09
`define CUBE_LUT_37AB 16'h2F0B
`define CUBE_LUT_37AC 16'h2F0E
`define CUBE_LUT_37AD 16'h2F11
`define CUBE_LUT_37AE 16'h2F14
`define CUBE_LUT_37AF 16'h2F16
`define CUBE_LUT_37B0 16'h2F19
`define CUBE_LUT_37B1 16'h2F1C
`define CUBE_LUT_37B2 16'h2F1F
`define CUBE_LUT_37B3 16'h2F22
`define CUBE_LUT_37B4 16'h2F24
`define CUBE_LUT_37B5 16'h2F27
`define CUBE_LUT_37B6 16'h2F2A
`define CUBE_LUT_37B7 16'h2F2D
`define CUBE_LUT_37B8 16'h2F30
`define CUBE_LUT_37B9 16'h2F32
`define CUBE_LUT_37BA 16'h2F35
`define CUBE_LUT_37BB 16'h2F38
`define CUBE_LUT_37BC 16'h2F3B
`define CUBE_LUT_37BD 16'h2F3E
`define CUBE_LUT_37BE 16'h2F40
`define CUBE_LUT_37BF 16'h2F43
`define CUBE_LUT_37C0 16'h2F46
`define CUBE_LUT_37C1 16'h2F49
`define CUBE_LUT_37C2 16'h2F4C
`define CUBE_LUT_37C3 16'h2F4E
`define CUBE_LUT_37C4 16'h2F51
`define CUBE_LUT_37C5 16'h2F54
`define CUBE_LUT_37C6 16'h2F57
`define CUBE_LUT_37C7 16'h2F5A
`define CUBE_LUT_37C8 16'h2F5D
`define CUBE_LUT_37C9 16'h2F5F
`define CUBE_LUT_37CA 16'h2F62
`define CUBE_LUT_37CB 16'h2F65
`define CUBE_LUT_37CC 16'h2F68
`define CUBE_LUT_37CD 16'h2F6B
`define CUBE_LUT_37CE 16'h2F6E
`define CUBE_LUT_37CF 16'h2F70
`define CUBE_LUT_37D0 16'h2F73
`define CUBE_LUT_37D1 16'h2F76
`define CUBE_LUT_37D2 16'h2F79
`define CUBE_LUT_37D3 16'h2F7C
`define CUBE_LUT_37D4 16'h2F7F
`define CUBE_LUT_37D5 16'h2F82
`define CUBE_LUT_37D6 16'h2F85
`define CUBE_LUT_37D7 16'h2F87
`define CUBE_LUT_37D8 16'h2F8A
`define CUBE_LUT_37D9 16'h2F8D
`define CUBE_LUT_37DA 16'h2F90
`define CUBE_LUT_37DB 16'h2F93
`define CUBE_LUT_37DC 16'h2F96
`define CUBE_LUT_37DD 16'h2F99
`define CUBE_LUT_37DE 16'h2F9C
`define CUBE_LUT_37DF 16'h2F9F
`define CUBE_LUT_37E0 16'h2FA1
`define CUBE_LUT_37E1 16'h2FA4
`define CUBE_LUT_37E2 16'h2FA7
`define CUBE_LUT_37E3 16'h2FAA
`define CUBE_LUT_37E4 16'h2FAD
`define CUBE_LUT_37E5 16'h2FB0
`define CUBE_LUT_37E6 16'h2FB3
`define CUBE_LUT_37E7 16'h2FB6
`define CUBE_LUT_37E8 16'h2FB9
`define CUBE_LUT_37E9 16'h2FBC
`define CUBE_LUT_37EA 16'h2FBF
`define CUBE_LUT_37EB 16'h2FC2
`define CUBE_LUT_37EC 16'h2FC5
`define CUBE_LUT_37ED 16'h2FC8
`define CUBE_LUT_37EE 16'h2FCA
`define CUBE_LUT_37EF 16'h2FCD
`define CUBE_LUT_37F0 16'h2FD0
`define CUBE_LUT_37F1 16'h2FD3
`define CUBE_LUT_37F2 16'h2FD6
`define CUBE_LUT_37F3 16'h2FD9
`define CUBE_LUT_37F4 16'h2FDC
`define CUBE_LUT_37F5 16'h2FDF
`define CUBE_LUT_37F6 16'h2FE2
`define CUBE_LUT_37F7 16'h2FE5
`define CUBE_LUT_37F8 16'h2FE8
`define CUBE_LUT_37F9 16'h2FEB
`define CUBE_LUT_37FA 16'h2FEE
`define CUBE_LUT_37FB 16'h2FF1
`define CUBE_LUT_37FC 16'h2FF4
`define CUBE_LUT_37FD 16'h2FF7
`define CUBE_LUT_37FE 16'h2FFA
`define CUBE_LUT_37FF 16'h2FFD
`define CUBE_LUT_3800 16'h3000
`define CUBE_LUT_3801 16'h3003
`define CUBE_LUT_3802 16'h3006
`define CUBE_LUT_3803 16'h3009
`define CUBE_LUT_3804 16'h300C
`define CUBE_LUT_3805 16'h300F
`define CUBE_LUT_3806 16'h3012
`define CUBE_LUT_3807 16'h3015
`define CUBE_LUT_3808 16'h3018
`define CUBE_LUT_3809 16'h301B
`define CUBE_LUT_380A 16'h301E
`define CUBE_LUT_380B 16'h3021
`define CUBE_LUT_380C 16'h3024
`define CUBE_LUT_380D 16'h3027
`define CUBE_LUT_380E 16'h302B
`define CUBE_LUT_380F 16'h302E
`define CUBE_LUT_3810 16'h3031
`define CUBE_LUT_3811 16'h3034
`define CUBE_LUT_3812 16'h3037
`define CUBE_LUT_3813 16'h303A
`define CUBE_LUT_3814 16'h303D
`define CUBE_LUT_3815 16'h3040
`define CUBE_LUT_3816 16'h3043
`define CUBE_LUT_3817 16'h3047
`define CUBE_LUT_3818 16'h304A
`define CUBE_LUT_3819 16'h304D
`define CUBE_LUT_381A 16'h3050
`define CUBE_LUT_381B 16'h3053
`define CUBE_LUT_381C 16'h3056
`define CUBE_LUT_381D 16'h3059
`define CUBE_LUT_381E 16'h305D
`define CUBE_LUT_381F 16'h3060
`define CUBE_LUT_3820 16'h3063
`define CUBE_LUT_3821 16'h3066
`define CUBE_LUT_3822 16'h3069
`define CUBE_LUT_3823 16'h306D
`define CUBE_LUT_3824 16'h3070
`define CUBE_LUT_3825 16'h3073
`define CUBE_LUT_3826 16'h3076
`define CUBE_LUT_3827 16'h307A
`define CUBE_LUT_3828 16'h307D
`define CUBE_LUT_3829 16'h3080
`define CUBE_LUT_382A 16'h3083
`define CUBE_LUT_382B 16'h3086
`define CUBE_LUT_382C 16'h308A
`define CUBE_LUT_382D 16'h308D
`define CUBE_LUT_382E 16'h3090
`define CUBE_LUT_382F 16'h3094
`define CUBE_LUT_3830 16'h3097
`define CUBE_LUT_3831 16'h309A
`define CUBE_LUT_3832 16'h309D
`define CUBE_LUT_3833 16'h30A1
`define CUBE_LUT_3834 16'h30A4
`define CUBE_LUT_3835 16'h30A7
`define CUBE_LUT_3836 16'h30AB
`define CUBE_LUT_3837 16'h30AE
`define CUBE_LUT_3838 16'h30B1
`define CUBE_LUT_3839 16'h30B5
`define CUBE_LUT_383A 16'h30B8
`define CUBE_LUT_383B 16'h30BB
`define CUBE_LUT_383C 16'h30BF
`define CUBE_LUT_383D 16'h30C2
`define CUBE_LUT_383E 16'h30C5
`define CUBE_LUT_383F 16'h30C9
`define CUBE_LUT_3840 16'h30CC
`define CUBE_LUT_3841 16'h30D0
`define CUBE_LUT_3842 16'h30D3
`define CUBE_LUT_3843 16'h30D6
`define CUBE_LUT_3844 16'h30DA
`define CUBE_LUT_3845 16'h30DD
`define CUBE_LUT_3846 16'h30E1
`define CUBE_LUT_3847 16'h30E4
`define CUBE_LUT_3848 16'h30E8
`define CUBE_LUT_3849 16'h30EB
`define CUBE_LUT_384A 16'h30EE
`define CUBE_LUT_384B 16'h30F2
`define CUBE_LUT_384C 16'h30F5
`define CUBE_LUT_384D 16'h30F9
`define CUBE_LUT_384E 16'h30FC
`define CUBE_LUT_384F 16'h3100
`define CUBE_LUT_3850 16'h3103
`define CUBE_LUT_3851 16'h3107
`define CUBE_LUT_3852 16'h310A
`define CUBE_LUT_3853 16'h310E
`define CUBE_LUT_3854 16'h3111
`define CUBE_LUT_3855 16'h3115
`define CUBE_LUT_3856 16'h3118
`define CUBE_LUT_3857 16'h311C
`define CUBE_LUT_3858 16'h311F
`define CUBE_LUT_3859 16'h3123
`define CUBE_LUT_385A 16'h3126
`define CUBE_LUT_385B 16'h312A
`define CUBE_LUT_385C 16'h312E
`define CUBE_LUT_385D 16'h3131
`define CUBE_LUT_385E 16'h3135
`define CUBE_LUT_385F 16'h3138
`define CUBE_LUT_3860 16'h313C
`define CUBE_LUT_3861 16'h313F
`define CUBE_LUT_3862 16'h3143
`define CUBE_LUT_3863 16'h3147
`define CUBE_LUT_3864 16'h314A
`define CUBE_LUT_3865 16'h314E
`define CUBE_LUT_3866 16'h3151
`define CUBE_LUT_3867 16'h3155
`define CUBE_LUT_3868 16'h3159
`define CUBE_LUT_3869 16'h315C
`define CUBE_LUT_386A 16'h3160
`define CUBE_LUT_386B 16'h3164
`define CUBE_LUT_386C 16'h3167
`define CUBE_LUT_386D 16'h316B
`define CUBE_LUT_386E 16'h316F
`define CUBE_LUT_386F 16'h3172
`define CUBE_LUT_3870 16'h3176
`define CUBE_LUT_3871 16'h317A
`define CUBE_LUT_3872 16'h317D
`define CUBE_LUT_3873 16'h3181
`define CUBE_LUT_3874 16'h3185
`define CUBE_LUT_3875 16'h3189
`define CUBE_LUT_3876 16'h318C
`define CUBE_LUT_3877 16'h3190
`define CUBE_LUT_3878 16'h3194
`define CUBE_LUT_3879 16'h3198
`define CUBE_LUT_387A 16'h319B
`define CUBE_LUT_387B 16'h319F
`define CUBE_LUT_387C 16'h31A3
`define CUBE_LUT_387D 16'h31A7
`define CUBE_LUT_387E 16'h31AA
`define CUBE_LUT_387F 16'h31AE
`define CUBE_LUT_3880 16'h31B2
`define CUBE_LUT_3881 16'h31B6
`define CUBE_LUT_3882 16'h31BA
`define CUBE_LUT_3883 16'h31BD
`define CUBE_LUT_3884 16'h31C1
`define CUBE_LUT_3885 16'h31C5
`define CUBE_LUT_3886 16'h31C9
`define CUBE_LUT_3887 16'h31CD
`define CUBE_LUT_3888 16'h31D1
`define CUBE_LUT_3889 16'h31D4
`define CUBE_LUT_388A 16'h31D8
`define CUBE_LUT_388B 16'h31DC
`define CUBE_LUT_388C 16'h31E0
`define CUBE_LUT_388D 16'h31E4
`define CUBE_LUT_388E 16'h31E8
`define CUBE_LUT_388F 16'h31EC
`define CUBE_LUT_3890 16'h31F0
`define CUBE_LUT_3891 16'h31F4
`define CUBE_LUT_3892 16'h31F7
`define CUBE_LUT_3893 16'h31FB
`define CUBE_LUT_3894 16'h31FF
`define CUBE_LUT_3895 16'h3203
`define CUBE_LUT_3896 16'h3207
`define CUBE_LUT_3897 16'h320B
`define CUBE_LUT_3898 16'h320F
`define CUBE_LUT_3899 16'h3213
`define CUBE_LUT_389A 16'h3217
`define CUBE_LUT_389B 16'h321B
`define CUBE_LUT_389C 16'h321F
`define CUBE_LUT_389D 16'h3223
`define CUBE_LUT_389E 16'h3227
`define CUBE_LUT_389F 16'h322B
`define CUBE_LUT_38A0 16'h322F
`define CUBE_LUT_38A1 16'h3233
`define CUBE_LUT_38A2 16'h3237
`define CUBE_LUT_38A3 16'h323B
`define CUBE_LUT_38A4 16'h323F
`define CUBE_LUT_38A5 16'h3243
`define CUBE_LUT_38A6 16'h3247
`define CUBE_LUT_38A7 16'h324B
`define CUBE_LUT_38A8 16'h324F
`define CUBE_LUT_38A9 16'h3253
`define CUBE_LUT_38AA 16'h3257
`define CUBE_LUT_38AB 16'h325B
`define CUBE_LUT_38AC 16'h3260
`define CUBE_LUT_38AD 16'h3264
`define CUBE_LUT_38AE 16'h3268
`define CUBE_LUT_38AF 16'h326C
`define CUBE_LUT_38B0 16'h3270
`define CUBE_LUT_38B1 16'h3274
`define CUBE_LUT_38B2 16'h3278
`define CUBE_LUT_38B3 16'h327C
`define CUBE_LUT_38B4 16'h3280
`define CUBE_LUT_38B5 16'h3285
`define CUBE_LUT_38B6 16'h3289
`define CUBE_LUT_38B7 16'h328D
`define CUBE_LUT_38B8 16'h3291
`define CUBE_LUT_38B9 16'h3295
`define CUBE_LUT_38BA 16'h3299
`define CUBE_LUT_38BB 16'h329E
`define CUBE_LUT_38BC 16'h32A2
`define CUBE_LUT_38BD 16'h32A6
`define CUBE_LUT_38BE 16'h32AA
`define CUBE_LUT_38BF 16'h32AF
`define CUBE_LUT_38C0 16'h32B3
`define CUBE_LUT_38C1 16'h32B7
`define CUBE_LUT_38C2 16'h32BB
`define CUBE_LUT_38C3 16'h32BF
`define CUBE_LUT_38C4 16'h32C4
`define CUBE_LUT_38C5 16'h32C8
`define CUBE_LUT_38C6 16'h32CC
`define CUBE_LUT_38C7 16'h32D1
`define CUBE_LUT_38C8 16'h32D5
`define CUBE_LUT_38C9 16'h32D9
`define CUBE_LUT_38CA 16'h32DD
`define CUBE_LUT_38CB 16'h32E2
`define CUBE_LUT_38CC 16'h32E6
`define CUBE_LUT_38CD 16'h32EA
`define CUBE_LUT_38CE 16'h32EF
`define CUBE_LUT_38CF 16'h32F3
`define CUBE_LUT_38D0 16'h32F7
`define CUBE_LUT_38D1 16'h32FC
`define CUBE_LUT_38D2 16'h3300
`define CUBE_LUT_38D3 16'h3304
`define CUBE_LUT_38D4 16'h3309
`define CUBE_LUT_38D5 16'h330D
`define CUBE_LUT_38D6 16'h3312
`define CUBE_LUT_38D7 16'h3316
`define CUBE_LUT_38D8 16'h331A
`define CUBE_LUT_38D9 16'h331F
`define CUBE_LUT_38DA 16'h3323
`define CUBE_LUT_38DB 16'h3328
`define CUBE_LUT_38DC 16'h332C
`define CUBE_LUT_38DD 16'h3330
`define CUBE_LUT_38DE 16'h3335
`define CUBE_LUT_38DF 16'h3339
`define CUBE_LUT_38E0 16'h333E
`define CUBE_LUT_38E1 16'h3342
`define CUBE_LUT_38E2 16'h3347
`define CUBE_LUT_38E3 16'h334B
`define CUBE_LUT_38E4 16'h3350
`define CUBE_LUT_38E5 16'h3354
`define CUBE_LUT_38E6 16'h3359
`define CUBE_LUT_38E7 16'h335D
`define CUBE_LUT_38E8 16'h3362
`define CUBE_LUT_38E9 16'h3366
`define CUBE_LUT_38EA 16'h336B
`define CUBE_LUT_38EB 16'h336F
`define CUBE_LUT_38EC 16'h3374
`define CUBE_LUT_38ED 16'h3378
`define CUBE_LUT_38EE 16'h337D
`define CUBE_LUT_38EF 16'h3381
`define CUBE_LUT_38F0 16'h3386
`define CUBE_LUT_38F1 16'h338B
`define CUBE_LUT_38F2 16'h338F
`define CUBE_LUT_38F3 16'h3394
`define CUBE_LUT_38F4 16'h3398
`define CUBE_LUT_38F5 16'h339D
`define CUBE_LUT_38F6 16'h33A1
`define CUBE_LUT_38F7 16'h33A6
`define CUBE_LUT_38F8 16'h33AB
`define CUBE_LUT_38F9 16'h33AF
`define CUBE_LUT_38FA 16'h33B4
`define CUBE_LUT_38FB 16'h33B9
`define CUBE_LUT_38FC 16'h33BD
`define CUBE_LUT_38FD 16'h33C2
`define CUBE_LUT_38FE 16'h33C7
`define CUBE_LUT_38FF 16'h33CB
`define CUBE_LUT_3900 16'h33D0
`define CUBE_LUT_3901 16'h33D5
`define CUBE_LUT_3902 16'h33D9
`define CUBE_LUT_3903 16'h33DE
`define CUBE_LUT_3904 16'h33E3
`define CUBE_LUT_3905 16'h33E8
`define CUBE_LUT_3906 16'h33EC
`define CUBE_LUT_3907 16'h33F1
`define CUBE_LUT_3908 16'h33F6
`define CUBE_LUT_3909 16'h33FA
`define CUBE_LUT_390A 16'h33FF
`define CUBE_LUT_390B 16'h3402
`define CUBE_LUT_390C 16'h3404
`define CUBE_LUT_390D 16'h3407
`define CUBE_LUT_390E 16'h3409
`define CUBE_LUT_390F 16'h340C
`define CUBE_LUT_3910 16'h340E
`define CUBE_LUT_3911 16'h3410
`define CUBE_LUT_3912 16'h3413
`define CUBE_LUT_3913 16'h3415
`define CUBE_LUT_3914 16'h3418
`define CUBE_LUT_3915 16'h341A
`define CUBE_LUT_3916 16'h341C
`define CUBE_LUT_3917 16'h341F
`define CUBE_LUT_3918 16'h3421
`define CUBE_LUT_3919 16'h3424
`define CUBE_LUT_391A 16'h3426
`define CUBE_LUT_391B 16'h3429
`define CUBE_LUT_391C 16'h342B
`define CUBE_LUT_391D 16'h342E
`define CUBE_LUT_391E 16'h3430
`define CUBE_LUT_391F 16'h3432
`define CUBE_LUT_3920 16'h3435
`define CUBE_LUT_3921 16'h3437
`define CUBE_LUT_3922 16'h343A
`define CUBE_LUT_3923 16'h343C
`define CUBE_LUT_3924 16'h343F
`define CUBE_LUT_3925 16'h3441
`define CUBE_LUT_3926 16'h3444
`define CUBE_LUT_3927 16'h3446
`define CUBE_LUT_3928 16'h3449
`define CUBE_LUT_3929 16'h344B
`define CUBE_LUT_392A 16'h344E
`define CUBE_LUT_392B 16'h3450
`define CUBE_LUT_392C 16'h3453
`define CUBE_LUT_392D 16'h3455
`define CUBE_LUT_392E 16'h3458
`define CUBE_LUT_392F 16'h345A
`define CUBE_LUT_3930 16'h345D
`define CUBE_LUT_3931 16'h345F
`define CUBE_LUT_3932 16'h3462
`define CUBE_LUT_3933 16'h3464
`define CUBE_LUT_3934 16'h3467
`define CUBE_LUT_3935 16'h3469
`define CUBE_LUT_3936 16'h346C
`define CUBE_LUT_3937 16'h346F
`define CUBE_LUT_3938 16'h3471
`define CUBE_LUT_3939 16'h3474
`define CUBE_LUT_393A 16'h3476
`define CUBE_LUT_393B 16'h3479
`define CUBE_LUT_393C 16'h347B
`define CUBE_LUT_393D 16'h347E
`define CUBE_LUT_393E 16'h3480
`define CUBE_LUT_393F 16'h3483
`define CUBE_LUT_3940 16'h3486
`define CUBE_LUT_3941 16'h3488
`define CUBE_LUT_3942 16'h348B
`define CUBE_LUT_3943 16'h348D
`define CUBE_LUT_3944 16'h3490
`define CUBE_LUT_3945 16'h3493
`define CUBE_LUT_3946 16'h3495
`define CUBE_LUT_3947 16'h3498
`define CUBE_LUT_3948 16'h349A
`define CUBE_LUT_3949 16'h349D
`define CUBE_LUT_394A 16'h34A0
`define CUBE_LUT_394B 16'h34A2
`define CUBE_LUT_394C 16'h34A5
`define CUBE_LUT_394D 16'h34A8
`define CUBE_LUT_394E 16'h34AA
`define CUBE_LUT_394F 16'h34AD
`define CUBE_LUT_3950 16'h34AF
`define CUBE_LUT_3951 16'h34B2
`define CUBE_LUT_3952 16'h34B5
`define CUBE_LUT_3953 16'h34B7
`define CUBE_LUT_3954 16'h34BA
`define CUBE_LUT_3955 16'h34BD
`define CUBE_LUT_3956 16'h34BF
`define CUBE_LUT_3957 16'h34C2
`define CUBE_LUT_3958 16'h34C5
`define CUBE_LUT_3959 16'h34C7
`define CUBE_LUT_395A 16'h34CA
`define CUBE_LUT_395B 16'h34CD
`define CUBE_LUT_395C 16'h34CF
`define CUBE_LUT_395D 16'h34D2
`define CUBE_LUT_395E 16'h34D5
`define CUBE_LUT_395F 16'h34D8
`define CUBE_LUT_3960 16'h34DA
`define CUBE_LUT_3961 16'h34DD
`define CUBE_LUT_3962 16'h34E0
`define CUBE_LUT_3963 16'h34E2
`define CUBE_LUT_3964 16'h34E5
`define CUBE_LUT_3965 16'h34E8
`define CUBE_LUT_3966 16'h34EB
`define CUBE_LUT_3967 16'h34ED
`define CUBE_LUT_3968 16'h34F0
`define CUBE_LUT_3969 16'h34F3
`define CUBE_LUT_396A 16'h34F6
`define CUBE_LUT_396B 16'h34F8
`define CUBE_LUT_396C 16'h34FB
`define CUBE_LUT_396D 16'h34FE
`define CUBE_LUT_396E 16'h3501
`define CUBE_LUT_396F 16'h3503
`define CUBE_LUT_3970 16'h3506
`define CUBE_LUT_3971 16'h3509
`define CUBE_LUT_3972 16'h350C
`define CUBE_LUT_3973 16'h350E
`define CUBE_LUT_3974 16'h3511
`define CUBE_LUT_3975 16'h3514
`define CUBE_LUT_3976 16'h3517
`define CUBE_LUT_3977 16'h351A
`define CUBE_LUT_3978 16'h351C
`define CUBE_LUT_3979 16'h351F
`define CUBE_LUT_397A 16'h3522
`define CUBE_LUT_397B 16'h3525
`define CUBE_LUT_397C 16'h3528
`define CUBE_LUT_397D 16'h352B
`define CUBE_LUT_397E 16'h352D
`define CUBE_LUT_397F 16'h3530
`define CUBE_LUT_3980 16'h3533
`define CUBE_LUT_3981 16'h3536
`define CUBE_LUT_3982 16'h3539
`define CUBE_LUT_3983 16'h353C
`define CUBE_LUT_3984 16'h353E
`define CUBE_LUT_3985 16'h3541
`define CUBE_LUT_3986 16'h3544
`define CUBE_LUT_3987 16'h3547
`define CUBE_LUT_3988 16'h354A
`define CUBE_LUT_3989 16'h354D
`define CUBE_LUT_398A 16'h3550
`define CUBE_LUT_398B 16'h3552
`define CUBE_LUT_398C 16'h3555
`define CUBE_LUT_398D 16'h3558
`define CUBE_LUT_398E 16'h355B
`define CUBE_LUT_398F 16'h355E
`define CUBE_LUT_3990 16'h3561
`define CUBE_LUT_3991 16'h3564
`define CUBE_LUT_3992 16'h3567
`define CUBE_LUT_3993 16'h356A
`define CUBE_LUT_3994 16'h356D
`define CUBE_LUT_3995 16'h356F
`define CUBE_LUT_3996 16'h3572
`define CUBE_LUT_3997 16'h3575
`define CUBE_LUT_3998 16'h3578
`define CUBE_LUT_3999 16'h357B
`define CUBE_LUT_399A 16'h357E
`define CUBE_LUT_399B 16'h3581
`define CUBE_LUT_399C 16'h3584
`define CUBE_LUT_399D 16'h3587
`define CUBE_LUT_399E 16'h358A
`define CUBE_LUT_399F 16'h358D
`define CUBE_LUT_39A0 16'h3590
`define CUBE_LUT_39A1 16'h3593
`define CUBE_LUT_39A2 16'h3596
`define CUBE_LUT_39A3 16'h3599
`define CUBE_LUT_39A4 16'h359C
`define CUBE_LUT_39A5 16'h359F
`define CUBE_LUT_39A6 16'h35A2
`define CUBE_LUT_39A7 16'h35A5
`define CUBE_LUT_39A8 16'h35A8
`define CUBE_LUT_39A9 16'h35AB
`define CUBE_LUT_39AA 16'h35AE
`define CUBE_LUT_39AB 16'h35B1
`define CUBE_LUT_39AC 16'h35B4
`define CUBE_LUT_39AD 16'h35B7
`define CUBE_LUT_39AE 16'h35BA
`define CUBE_LUT_39AF 16'h35BD
`define CUBE_LUT_39B0 16'h35C0
`define CUBE_LUT_39B1 16'h35C3
`define CUBE_LUT_39B2 16'h35C6
`define CUBE_LUT_39B3 16'h35C9
`define CUBE_LUT_39B4 16'h35CC
`define CUBE_LUT_39B5 16'h35CF
`define CUBE_LUT_39B6 16'h35D2
`define CUBE_LUT_39B7 16'h35D5
`define CUBE_LUT_39B8 16'h35D8
`define CUBE_LUT_39B9 16'h35DB
`define CUBE_LUT_39BA 16'h35DE
`define CUBE_LUT_39BB 16'h35E1
`define CUBE_LUT_39BC 16'h35E5
`define CUBE_LUT_39BD 16'h35E8
`define CUBE_LUT_39BE 16'h35EB
`define CUBE_LUT_39BF 16'h35EE
`define CUBE_LUT_39C0 16'h35F1
`define CUBE_LUT_39C1 16'h35F4
`define CUBE_LUT_39C2 16'h35F7
`define CUBE_LUT_39C3 16'h35FA
`define CUBE_LUT_39C4 16'h35FD
`define CUBE_LUT_39C5 16'h3600
`define CUBE_LUT_39C6 16'h3604
`define CUBE_LUT_39C7 16'h3607
`define CUBE_LUT_39C8 16'h360A
`define CUBE_LUT_39C9 16'h360D
`define CUBE_LUT_39CA 16'h3610
`define CUBE_LUT_39CB 16'h3613
`define CUBE_LUT_39CC 16'h3616
`define CUBE_LUT_39CD 16'h361A
`define CUBE_LUT_39CE 16'h361D
`define CUBE_LUT_39CF 16'h3620
`define CUBE_LUT_39D0 16'h3623
`define CUBE_LUT_39D1 16'h3626
`define CUBE_LUT_39D2 16'h3629
`define CUBE_LUT_39D3 16'h362D
`define CUBE_LUT_39D4 16'h3630
`define CUBE_LUT_39D5 16'h3633
`define CUBE_LUT_39D6 16'h3636
`define CUBE_LUT_39D7 16'h3639
`define CUBE_LUT_39D8 16'h363C
`define CUBE_LUT_39D9 16'h3640
`define CUBE_LUT_39DA 16'h3643
`define CUBE_LUT_39DB 16'h3646
`define CUBE_LUT_39DC 16'h3649
`define CUBE_LUT_39DD 16'h364D
`define CUBE_LUT_39DE 16'h3650
`define CUBE_LUT_39DF 16'h3653
`define CUBE_LUT_39E0 16'h3656
`define CUBE_LUT_39E1 16'h3659
`define CUBE_LUT_39E2 16'h365D
`define CUBE_LUT_39E3 16'h3660
`define CUBE_LUT_39E4 16'h3663
`define CUBE_LUT_39E5 16'h3666
`define CUBE_LUT_39E6 16'h366A
`define CUBE_LUT_39E7 16'h366D
`define CUBE_LUT_39E8 16'h3670
`define CUBE_LUT_39E9 16'h3674
`define CUBE_LUT_39EA 16'h3677
`define CUBE_LUT_39EB 16'h367A
`define CUBE_LUT_39EC 16'h367D
`define CUBE_LUT_39ED 16'h3681
`define CUBE_LUT_39EE 16'h3684
`define CUBE_LUT_39EF 16'h3687
`define CUBE_LUT_39F0 16'h368B
`define CUBE_LUT_39F1 16'h368E
`define CUBE_LUT_39F2 16'h3691
`define CUBE_LUT_39F3 16'h3694
`define CUBE_LUT_39F4 16'h3698
`define CUBE_LUT_39F5 16'h369B
`define CUBE_LUT_39F6 16'h369E
`define CUBE_LUT_39F7 16'h36A2
`define CUBE_LUT_39F8 16'h36A5
`define CUBE_LUT_39F9 16'h36A8
`define CUBE_LUT_39FA 16'h36AC
`define CUBE_LUT_39FB 16'h36AF
`define CUBE_LUT_39FC 16'h36B3
`define CUBE_LUT_39FD 16'h36B6
`define CUBE_LUT_39FE 16'h36B9
`define CUBE_LUT_39FF 16'h36BD
`define CUBE_LUT_3A00 16'h36C0
`define CUBE_LUT_3A01 16'h36C3
`define CUBE_LUT_3A02 16'h36C7
`define CUBE_LUT_3A03 16'h36CA
`define CUBE_LUT_3A04 16'h36CE
`define CUBE_LUT_3A05 16'h36D1
`define CUBE_LUT_3A06 16'h36D4
`define CUBE_LUT_3A07 16'h36D8
`define CUBE_LUT_3A08 16'h36DB
`define CUBE_LUT_3A09 16'h36DF
`define CUBE_LUT_3A0A 16'h36E2
`define CUBE_LUT_3A0B 16'h36E5
`define CUBE_LUT_3A0C 16'h36E9
`define CUBE_LUT_3A0D 16'h36EC
`define CUBE_LUT_3A0E 16'h36F0
`define CUBE_LUT_3A0F 16'h36F3
`define CUBE_LUT_3A10 16'h36F7
`define CUBE_LUT_3A11 16'h36FA
`define CUBE_LUT_3A12 16'h36FD
`define CUBE_LUT_3A13 16'h3701
`define CUBE_LUT_3A14 16'h3704
`define CUBE_LUT_3A15 16'h3708
`define CUBE_LUT_3A16 16'h370B
`define CUBE_LUT_3A17 16'h370F
`define CUBE_LUT_3A18 16'h3712
`define CUBE_LUT_3A19 16'h3716
`define CUBE_LUT_3A1A 16'h3719
`define CUBE_LUT_3A1B 16'h371D
`define CUBE_LUT_3A1C 16'h3720
`define CUBE_LUT_3A1D 16'h3724
`define CUBE_LUT_3A1E 16'h3727
`define CUBE_LUT_3A1F 16'h372B
`define CUBE_LUT_3A20 16'h372E
`define CUBE_LUT_3A21 16'h3732
`define CUBE_LUT_3A22 16'h3735
`define CUBE_LUT_3A23 16'h3739
`define CUBE_LUT_3A24 16'h373C
`define CUBE_LUT_3A25 16'h3740
`define CUBE_LUT_3A26 16'h3743
`define CUBE_LUT_3A27 16'h3747
`define CUBE_LUT_3A28 16'h374B
`define CUBE_LUT_3A29 16'h374E
`define CUBE_LUT_3A2A 16'h3752
`define CUBE_LUT_3A2B 16'h3755
`define CUBE_LUT_3A2C 16'h3759
`define CUBE_LUT_3A2D 16'h375C
`define CUBE_LUT_3A2E 16'h3760
`define CUBE_LUT_3A2F 16'h3764
`define CUBE_LUT_3A30 16'h3767
`define CUBE_LUT_3A31 16'h376B
`define CUBE_LUT_3A32 16'h376E
`define CUBE_LUT_3A33 16'h3772
`define CUBE_LUT_3A34 16'h3776
`define CUBE_LUT_3A35 16'h3779
`define CUBE_LUT_3A36 16'h377D
`define CUBE_LUT_3A37 16'h3780
`define CUBE_LUT_3A38 16'h3784
`define CUBE_LUT_3A39 16'h3788
`define CUBE_LUT_3A3A 16'h378B
`define CUBE_LUT_3A3B 16'h378F
`define CUBE_LUT_3A3C 16'h3793
`define CUBE_LUT_3A3D 16'h3796
`define CUBE_LUT_3A3E 16'h379A
`define CUBE_LUT_3A3F 16'h379D
`define CUBE_LUT_3A40 16'h37A1
`define CUBE_LUT_3A41 16'h37A5
`define CUBE_LUT_3A42 16'h37A8
`define CUBE_LUT_3A43 16'h37AC
`define CUBE_LUT_3A44 16'h37B0
`define CUBE_LUT_3A45 16'h37B3
`define CUBE_LUT_3A46 16'h37B7
`define CUBE_LUT_3A47 16'h37BB
`define CUBE_LUT_3A48 16'h37BF
`define CUBE_LUT_3A49 16'h37C2
`define CUBE_LUT_3A4A 16'h37C6
`define CUBE_LUT_3A4B 16'h37CA
`define CUBE_LUT_3A4C 16'h37CD
`define CUBE_LUT_3A4D 16'h37D1
`define CUBE_LUT_3A4E 16'h37D5
`define CUBE_LUT_3A4F 16'h37D9
`define CUBE_LUT_3A50 16'h37DC
`define CUBE_LUT_3A51 16'h37E0
`define CUBE_LUT_3A52 16'h37E4
`define CUBE_LUT_3A53 16'h37E8
`define CUBE_LUT_3A54 16'h37EB
`define CUBE_LUT_3A55 16'h37EF
`define CUBE_LUT_3A56 16'h37F3
`define CUBE_LUT_3A57 16'h37F7
`define CUBE_LUT_3A58 16'h37FA
`define CUBE_LUT_3A59 16'h37FE
`define CUBE_LUT_3A5A 16'h3801
`define CUBE_LUT_3A5B 16'h3803
`define CUBE_LUT_3A5C 16'h3805
`define CUBE_LUT_3A5D 16'h3807
`define CUBE_LUT_3A5E 16'h3809
`define CUBE_LUT_3A5F 16'h380A
`define CUBE_LUT_3A60 16'h380C
`define CUBE_LUT_3A61 16'h380E
`define CUBE_LUT_3A62 16'h3810
`define CUBE_LUT_3A63 16'h3812
`define CUBE_LUT_3A64 16'h3814
`define CUBE_LUT_3A65 16'h3816
`define CUBE_LUT_3A66 16'h3818
`define CUBE_LUT_3A67 16'h381A
`define CUBE_LUT_3A68 16'h381C
`define CUBE_LUT_3A69 16'h381E
`define CUBE_LUT_3A6A 16'h3820
`define CUBE_LUT_3A6B 16'h3821
`define CUBE_LUT_3A6C 16'h3823
`define CUBE_LUT_3A6D 16'h3825
`define CUBE_LUT_3A6E 16'h3827
`define CUBE_LUT_3A6F 16'h3829
`define CUBE_LUT_3A70 16'h382B
`define CUBE_LUT_3A71 16'h382D
`define CUBE_LUT_3A72 16'h382F
`define CUBE_LUT_3A73 16'h3831
`define CUBE_LUT_3A74 16'h3833
`define CUBE_LUT_3A75 16'h3835
`define CUBE_LUT_3A76 16'h3837
`define CUBE_LUT_3A77 16'h3839
`define CUBE_LUT_3A78 16'h383B
`define CUBE_LUT_3A79 16'h383D
`define CUBE_LUT_3A7A 16'h383F
`define CUBE_LUT_3A7B 16'h3841
`define CUBE_LUT_3A7C 16'h3843
`define CUBE_LUT_3A7D 16'h3845
`define CUBE_LUT_3A7E 16'h3847
`define CUBE_LUT_3A7F 16'h3849
`define CUBE_LUT_3A80 16'h384A
`define CUBE_LUT_3A81 16'h384C
`define CUBE_LUT_3A82 16'h384E
`define CUBE_LUT_3A83 16'h3850
`define CUBE_LUT_3A84 16'h3852
`define CUBE_LUT_3A85 16'h3854
`define CUBE_LUT_3A86 16'h3856
`define CUBE_LUT_3A87 16'h3858
`define CUBE_LUT_3A88 16'h385A
`define CUBE_LUT_3A89 16'h385C
`define CUBE_LUT_3A8A 16'h385E
`define CUBE_LUT_3A8B 16'h3860
`define CUBE_LUT_3A8C 16'h3862
`define CUBE_LUT_3A8D 16'h3864
`define CUBE_LUT_3A8E 16'h3866
`define CUBE_LUT_3A8F 16'h3868
`define CUBE_LUT_3A90 16'h386A
`define CUBE_LUT_3A91 16'h386D
`define CUBE_LUT_3A92 16'h386F
`define CUBE_LUT_3A93 16'h3871
`define CUBE_LUT_3A94 16'h3873
`define CUBE_LUT_3A95 16'h3875
`define CUBE_LUT_3A96 16'h3877
`define CUBE_LUT_3A97 16'h3879
`define CUBE_LUT_3A98 16'h387B
`define CUBE_LUT_3A99 16'h387D
`define CUBE_LUT_3A9A 16'h387F
`define CUBE_LUT_3A9B 16'h3881
`define CUBE_LUT_3A9C 16'h3883
`define CUBE_LUT_3A9D 16'h3885
`define CUBE_LUT_3A9E 16'h3887
`define CUBE_LUT_3A9F 16'h3889
`define CUBE_LUT_3AA0 16'h388B
`define CUBE_LUT_3AA1 16'h388D
`define CUBE_LUT_3AA2 16'h388F
`define CUBE_LUT_3AA3 16'h3891
`define CUBE_LUT_3AA4 16'h3893
`define CUBE_LUT_3AA5 16'h3895
`define CUBE_LUT_3AA6 16'h3897
`define CUBE_LUT_3AA7 16'h389A
`define CUBE_LUT_3AA8 16'h389C
`define CUBE_LUT_3AA9 16'h389E
`define CUBE_LUT_3AAA 16'h38A0
`define CUBE_LUT_3AAB 16'h38A2
`define CUBE_LUT_3AAC 16'h38A4
`define CUBE_LUT_3AAD 16'h38A6
`define CUBE_LUT_3AAE 16'h38A8
`define CUBE_LUT_3AAF 16'h38AA
`define CUBE_LUT_3AB0 16'h38AC
`define CUBE_LUT_3AB1 16'h38AE
`define CUBE_LUT_3AB2 16'h38B1
`define CUBE_LUT_3AB3 16'h38B3
`define CUBE_LUT_3AB4 16'h38B5
`define CUBE_LUT_3AB5 16'h38B7
`define CUBE_LUT_3AB6 16'h38B9
`define CUBE_LUT_3AB7 16'h38BB
`define CUBE_LUT_3AB8 16'h38BD
`define CUBE_LUT_3AB9 16'h38BF
`define CUBE_LUT_3ABA 16'h38C1
`define CUBE_LUT_3ABB 16'h38C4
`define CUBE_LUT_3ABC 16'h38C6
`define CUBE_LUT_3ABD 16'h38C8
`define CUBE_LUT_3ABE 16'h38CA
`define CUBE_LUT_3ABF 16'h38CC
`define CUBE_LUT_3AC0 16'h38CE
`define CUBE_LUT_3AC1 16'h38D0
`define CUBE_LUT_3AC2 16'h38D2
`define CUBE_LUT_3AC3 16'h38D5
`define CUBE_LUT_3AC4 16'h38D7
`define CUBE_LUT_3AC5 16'h38D9
`define CUBE_LUT_3AC6 16'h38DB
`define CUBE_LUT_3AC7 16'h38DD
`define CUBE_LUT_3AC8 16'h38DF
`define CUBE_LUT_3AC9 16'h38E2
`define CUBE_LUT_3ACA 16'h38E4
`define CUBE_LUT_3ACB 16'h38E6
`define CUBE_LUT_3ACC 16'h38E8
`define CUBE_LUT_3ACD 16'h38EA
`define CUBE_LUT_3ACE 16'h38EC
`define CUBE_LUT_3ACF 16'h38EF
`define CUBE_LUT_3AD0 16'h38F1
`define CUBE_LUT_3AD1 16'h38F3
`define CUBE_LUT_3AD2 16'h38F5
`define CUBE_LUT_3AD3 16'h38F7
`define CUBE_LUT_3AD4 16'h38F9
`define CUBE_LUT_3AD5 16'h38FC
`define CUBE_LUT_3AD6 16'h38FE
`define CUBE_LUT_3AD7 16'h3900
`define CUBE_LUT_3AD8 16'h3902
`define CUBE_LUT_3AD9 16'h3904
`define CUBE_LUT_3ADA 16'h3907
`define CUBE_LUT_3ADB 16'h3909
`define CUBE_LUT_3ADC 16'h390B
`define CUBE_LUT_3ADD 16'h390D
`define CUBE_LUT_3ADE 16'h390F
`define CUBE_LUT_3ADF 16'h3912
`define CUBE_LUT_3AE0 16'h3914
`define CUBE_LUT_3AE1 16'h3916
`define CUBE_LUT_3AE2 16'h3918
`define CUBE_LUT_3AE3 16'h391A
`define CUBE_LUT_3AE4 16'h391D
`define CUBE_LUT_3AE5 16'h391F
`define CUBE_LUT_3AE6 16'h3921
`define CUBE_LUT_3AE7 16'h3923
`define CUBE_LUT_3AE8 16'h3926
`define CUBE_LUT_3AE9 16'h3928
`define CUBE_LUT_3AEA 16'h392A
`define CUBE_LUT_3AEB 16'h392C
`define CUBE_LUT_3AEC 16'h392F
`define CUBE_LUT_3AED 16'h3931
`define CUBE_LUT_3AEE 16'h3933
`define CUBE_LUT_3AEF 16'h3935
`define CUBE_LUT_3AF0 16'h3938
`define CUBE_LUT_3AF1 16'h393A
`define CUBE_LUT_3AF2 16'h393C
`define CUBE_LUT_3AF3 16'h393E
`define CUBE_LUT_3AF4 16'h3941
`define CUBE_LUT_3AF5 16'h3943
`define CUBE_LUT_3AF6 16'h3945
`define CUBE_LUT_3AF7 16'h3947
`define CUBE_LUT_3AF8 16'h394A
`define CUBE_LUT_3AF9 16'h394C
`define CUBE_LUT_3AFA 16'h394E
`define CUBE_LUT_3AFB 16'h3951
`define CUBE_LUT_3AFC 16'h3953
`define CUBE_LUT_3AFD 16'h3955
`define CUBE_LUT_3AFE 16'h3957
`define CUBE_LUT_3AFF 16'h395A
`define CUBE_LUT_3B00 16'h395C
`define CUBE_LUT_3B01 16'h395E
`define CUBE_LUT_3B02 16'h3961
`define CUBE_LUT_3B03 16'h3963
`define CUBE_LUT_3B04 16'h3965
`define CUBE_LUT_3B05 16'h3968
`define CUBE_LUT_3B06 16'h396A
`define CUBE_LUT_3B07 16'h396C
`define CUBE_LUT_3B08 16'h396E
`define CUBE_LUT_3B09 16'h3971
`define CUBE_LUT_3B0A 16'h3973
`define CUBE_LUT_3B0B 16'h3975
`define CUBE_LUT_3B0C 16'h3978
`define CUBE_LUT_3B0D 16'h397A
`define CUBE_LUT_3B0E 16'h397C
`define CUBE_LUT_3B0F 16'h397F
`define CUBE_LUT_3B10 16'h3981
`define CUBE_LUT_3B11 16'h3983
`define CUBE_LUT_3B12 16'h3986
`define CUBE_LUT_3B13 16'h3988
`define CUBE_LUT_3B14 16'h398A
`define CUBE_LUT_3B15 16'h398D
`define CUBE_LUT_3B16 16'h398F
`define CUBE_LUT_3B17 16'h3992
`define CUBE_LUT_3B18 16'h3994
`define CUBE_LUT_3B19 16'h3996
`define CUBE_LUT_3B1A 16'h3999
`define CUBE_LUT_3B1B 16'h399B
`define CUBE_LUT_3B1C 16'h399D
`define CUBE_LUT_3B1D 16'h39A0
`define CUBE_LUT_3B1E 16'h39A2
`define CUBE_LUT_3B1F 16'h39A4
`define CUBE_LUT_3B20 16'h39A7
`define CUBE_LUT_3B21 16'h39A9
`define CUBE_LUT_3B22 16'h39AC
`define CUBE_LUT_3B23 16'h39AE
`define CUBE_LUT_3B24 16'h39B0
`define CUBE_LUT_3B25 16'h39B3
`define CUBE_LUT_3B26 16'h39B5
`define CUBE_LUT_3B27 16'h39B8
`define CUBE_LUT_3B28 16'h39BA
`define CUBE_LUT_3B29 16'h39BC
`define CUBE_LUT_3B2A 16'h39BF
`define CUBE_LUT_3B2B 16'h39C1
`define CUBE_LUT_3B2C 16'h39C4
`define CUBE_LUT_3B2D 16'h39C6
`define CUBE_LUT_3B2E 16'h39C8
`define CUBE_LUT_3B2F 16'h39CB
`define CUBE_LUT_3B30 16'h39CD
`define CUBE_LUT_3B31 16'h39D0
`define CUBE_LUT_3B32 16'h39D2
`define CUBE_LUT_3B33 16'h39D5
`define CUBE_LUT_3B34 16'h39D7
`define CUBE_LUT_3B35 16'h39D9
`define CUBE_LUT_3B36 16'h39DC
`define CUBE_LUT_3B37 16'h39DE
`define CUBE_LUT_3B38 16'h39E1
`define CUBE_LUT_3B39 16'h39E3
`define CUBE_LUT_3B3A 16'h39E6
`define CUBE_LUT_3B3B 16'h39E8
`define CUBE_LUT_3B3C 16'h39EA
`define CUBE_LUT_3B3D 16'h39ED
`define CUBE_LUT_3B3E 16'h39EF
`define CUBE_LUT_3B3F 16'h39F2
`define CUBE_LUT_3B40 16'h39F4
`define CUBE_LUT_3B41 16'h39F7
`define CUBE_LUT_3B42 16'h39F9
`define CUBE_LUT_3B43 16'h39FC
`define CUBE_LUT_3B44 16'h39FE
`define CUBE_LUT_3B45 16'h3A01
`define CUBE_LUT_3B46 16'h3A03
`define CUBE_LUT_3B47 16'h3A06
`define CUBE_LUT_3B48 16'h3A08
`define CUBE_LUT_3B49 16'h3A0B
`define CUBE_LUT_3B4A 16'h3A0D
`define CUBE_LUT_3B4B 16'h3A10
`define CUBE_LUT_3B4C 16'h3A12
`define CUBE_LUT_3B4D 16'h3A15
`define CUBE_LUT_3B4E 16'h3A17
`define CUBE_LUT_3B4F 16'h3A1A
`define CUBE_LUT_3B50 16'h3A1C
`define CUBE_LUT_3B51 16'h3A1F
`define CUBE_LUT_3B52 16'h3A21
`define CUBE_LUT_3B53 16'h3A24
`define CUBE_LUT_3B54 16'h3A26
`define CUBE_LUT_3B55 16'h3A29
`define CUBE_LUT_3B56 16'h3A2B
`define CUBE_LUT_3B57 16'h3A2E
`define CUBE_LUT_3B58 16'h3A30
`define CUBE_LUT_3B59 16'h3A33
`define CUBE_LUT_3B5A 16'h3A35
`define CUBE_LUT_3B5B 16'h3A38
`define CUBE_LUT_3B5C 16'h3A3A
`define CUBE_LUT_3B5D 16'h3A3D
`define CUBE_LUT_3B5E 16'h3A3F
`define CUBE_LUT_3B5F 16'h3A42
`define CUBE_LUT_3B60 16'h3A45
`define CUBE_LUT_3B61 16'h3A47
`define CUBE_LUT_3B62 16'h3A4A
`define CUBE_LUT_3B63 16'h3A4C
`define CUBE_LUT_3B64 16'h3A4F
`define CUBE_LUT_3B65 16'h3A51
`define CUBE_LUT_3B66 16'h3A54
`define CUBE_LUT_3B67 16'h3A56
`define CUBE_LUT_3B68 16'h3A59
`define CUBE_LUT_3B69 16'h3A5C
`define CUBE_LUT_3B6A 16'h3A5E
`define CUBE_LUT_3B6B 16'h3A61
`define CUBE_LUT_3B6C 16'h3A63
`define CUBE_LUT_3B6D 16'h3A66
`define CUBE_LUT_3B6E 16'h3A68
`define CUBE_LUT_3B6F 16'h3A6B
`define CUBE_LUT_3B70 16'h3A6E
`define CUBE_LUT_3B71 16'h3A70
`define CUBE_LUT_3B72 16'h3A73
`define CUBE_LUT_3B73 16'h3A75
`define CUBE_LUT_3B74 16'h3A78
`define CUBE_LUT_3B75 16'h3A7B
`define CUBE_LUT_3B76 16'h3A7D
`define CUBE_LUT_3B77 16'h3A80
`define CUBE_LUT_3B78 16'h3A82
`define CUBE_LUT_3B79 16'h3A85
`define CUBE_LUT_3B7A 16'h3A88
`define CUBE_LUT_3B7B 16'h3A8A
`define CUBE_LUT_3B7C 16'h3A8D
`define CUBE_LUT_3B7D 16'h3A90
`define CUBE_LUT_3B7E 16'h3A92
`define CUBE_LUT_3B7F 16'h3A95
`define CUBE_LUT_3B80 16'h3A98
`define CUBE_LUT_3B81 16'h3A9A
`define CUBE_LUT_3B82 16'h3A9D
`define CUBE_LUT_3B83 16'h3A9F
`define CUBE_LUT_3B84 16'h3AA2
`define CUBE_LUT_3B85 16'h3AA5
`define CUBE_LUT_3B86 16'h3AA7
`define CUBE_LUT_3B87 16'h3AAA
`define CUBE_LUT_3B88 16'h3AAD
`define CUBE_LUT_3B89 16'h3AAF
`define CUBE_LUT_3B8A 16'h3AB2
`define CUBE_LUT_3B8B 16'h3AB5
`define CUBE_LUT_3B8C 16'h3AB7
`define CUBE_LUT_3B8D 16'h3ABA
`define CUBE_LUT_3B8E 16'h3ABD
`define CUBE_LUT_3B8F 16'h3ABF
`define CUBE_LUT_3B90 16'h3AC2
`define CUBE_LUT_3B91 16'h3AC5
`define CUBE_LUT_3B92 16'h3AC7
`define CUBE_LUT_3B93 16'h3ACA
`define CUBE_LUT_3B94 16'h3ACD
`define CUBE_LUT_3B95 16'h3ACF
`define CUBE_LUT_3B96 16'h3AD2
`define CUBE_LUT_3B97 16'h3AD5
`define CUBE_LUT_3B98 16'h3AD8
`define CUBE_LUT_3B99 16'h3ADA
`define CUBE_LUT_3B9A 16'h3ADD
`define CUBE_LUT_3B9B 16'h3AE0
`define CUBE_LUT_3B9C 16'h3AE2
`define CUBE_LUT_3B9D 16'h3AE5
`define CUBE_LUT_3B9E 16'h3AE8
`define CUBE_LUT_3B9F 16'h3AEB
`define CUBE_LUT_3BA0 16'h3AED
`define CUBE_LUT_3BA1 16'h3AF0
`define CUBE_LUT_3BA2 16'h3AF3
`define CUBE_LUT_3BA3 16'h3AF5
`define CUBE_LUT_3BA4 16'h3AF8
`define CUBE_LUT_3BA5 16'h3AFB
`define CUBE_LUT_3BA6 16'h3AFE
`define CUBE_LUT_3BA7 16'h3B00
`define CUBE_LUT_3BA8 16'h3B03
`define CUBE_LUT_3BA9 16'h3B06
`define CUBE_LUT_3BAA 16'h3B09
`define CUBE_LUT_3BAB 16'h3B0B
`define CUBE_LUT_3BAC 16'h3B0E
`define CUBE_LUT_3BAD 16'h3B11
`define CUBE_LUT_3BAE 16'h3B14
`define CUBE_LUT_3BAF 16'h3B16
`define CUBE_LUT_3BB0 16'h3B19
`define CUBE_LUT_3BB1 16'h3B1C
`define CUBE_LUT_3BB2 16'h3B1F
`define CUBE_LUT_3BB3 16'h3B22
`define CUBE_LUT_3BB4 16'h3B24
`define CUBE_LUT_3BB5 16'h3B27
`define CUBE_LUT_3BB6 16'h3B2A
`define CUBE_LUT_3BB7 16'h3B2D
`define CUBE_LUT_3BB8 16'h3B30
`define CUBE_LUT_3BB9 16'h3B32
`define CUBE_LUT_3BBA 16'h3B35
`define CUBE_LUT_3BBB 16'h3B38
`define CUBE_LUT_3BBC 16'h3B3B
`define CUBE_LUT_3BBD 16'h3B3E
`define CUBE_LUT_3BBE 16'h3B40
`define CUBE_LUT_3BBF 16'h3B43
`define CUBE_LUT_3BC0 16'h3B46
`define CUBE_LUT_3BC1 16'h3B49
`define CUBE_LUT_3BC2 16'h3B4C
`define CUBE_LUT_3BC3 16'h3B4E
`define CUBE_LUT_3BC4 16'h3B51
`define CUBE_LUT_3BC5 16'h3B54
`define CUBE_LUT_3BC6 16'h3B57
`define CUBE_LUT_3BC7 16'h3B5A
`define CUBE_LUT_3BC8 16'h3B5D
`define CUBE_LUT_3BC9 16'h3B5F
`define CUBE_LUT_3BCA 16'h3B62
`define CUBE_LUT_3BCB 16'h3B65
`define CUBE_LUT_3BCC 16'h3B68
`define CUBE_LUT_3BCD 16'h3B6B
`define CUBE_LUT_3BCE 16'h3B6E
`define CUBE_LUT_3BCF 16'h3B70
`define CUBE_LUT_3BD0 16'h3B73
`define CUBE_LUT_3BD1 16'h3B76
`define CUBE_LUT_3BD2 16'h3B79
`define CUBE_LUT_3BD3 16'h3B7C
`define CUBE_LUT_3BD4 16'h3B7F
`define CUBE_LUT_3BD5 16'h3B82
`define CUBE_LUT_3BD6 16'h3B85
`define CUBE_LUT_3BD7 16'h3B87
`define CUBE_LUT_3BD8 16'h3B8A
`define CUBE_LUT_3BD9 16'h3B8D
`define CUBE_LUT_3BDA 16'h3B90
`define CUBE_LUT_3BDB 16'h3B93
`define CUBE_LUT_3BDC 16'h3B96
`define CUBE_LUT_3BDD 16'h3B99
`define CUBE_LUT_3BDE 16'h3B9C
`define CUBE_LUT_3BDF 16'h3B9F
`define CUBE_LUT_3BE0 16'h3BA1
`define CUBE_LUT_3BE1 16'h3BA4
`define CUBE_LUT_3BE2 16'h3BA7
`define CUBE_LUT_3BE3 16'h3BAA
`define CUBE_LUT_3BE4 16'h3BAD
`define CUBE_LUT_3BE5 16'h3BB0
`define CUBE_LUT_3BE6 16'h3BB3
`define CUBE_LUT_3BE7 16'h3BB6
`define CUBE_LUT_3BE8 16'h3BB9
`define CUBE_LUT_3BE9 16'h3BBC
`define CUBE_LUT_3BEA 16'h3BBF
`define CUBE_LUT_3BEB 16'h3BC2
`define CUBE_LUT_3BEC 16'h3BC5
`define CUBE_LUT_3BED 16'h3BC8
`define CUBE_LUT_3BEE 16'h3BCA
`define CUBE_LUT_3BEF 16'h3BCD
`define CUBE_LUT_3BF0 16'h3BD0
`define CUBE_LUT_3BF1 16'h3BD3
`define CUBE_LUT_3BF2 16'h3BD6
`define CUBE_LUT_3BF3 16'h3BD9
`define CUBE_LUT_3BF4 16'h3BDC
`define CUBE_LUT_3BF5 16'h3BDF
`define CUBE_LUT_3BF6 16'h3BE2
`define CUBE_LUT_3BF7 16'h3BE5
`define CUBE_LUT_3BF8 16'h3BE8
`define CUBE_LUT_3BF9 16'h3BEB
`define CUBE_LUT_3BFA 16'h3BEE
`define CUBE_LUT_3BFB 16'h3BF1
`define CUBE_LUT_3BFC 16'h3BF4
`define CUBE_LUT_3BFD 16'h3BF7
`define CUBE_LUT_3BFE 16'h3BFA
`define CUBE_LUT_3BFF 16'h3BFD
`define CUBE_LUT_3C00 16'h3C00
`define CUBE_LUT_3C01 16'h3C03
`define CUBE_LUT_3C02 16'h3C06
`define CUBE_LUT_3C03 16'h3C09
`define CUBE_LUT_3C04 16'h3C0C
`define CUBE_LUT_3C05 16'h3C0F
`define CUBE_LUT_3C06 16'h3C12
`define CUBE_LUT_3C07 16'h3C15
`define CUBE_LUT_3C08 16'h3C18
`define CUBE_LUT_3C09 16'h3C1B
`define CUBE_LUT_3C0A 16'h3C1E
`define CUBE_LUT_3C0B 16'h3C21
`define CUBE_LUT_3C0C 16'h3C24
`define CUBE_LUT_3C0D 16'h3C27
`define CUBE_LUT_3C0E 16'h3C2B
`define CUBE_LUT_3C0F 16'h3C2E
`define CUBE_LUT_3C10 16'h3C31
`define CUBE_LUT_3C11 16'h3C34
`define CUBE_LUT_3C12 16'h3C37
`define CUBE_LUT_3C13 16'h3C3A
`define CUBE_LUT_3C14 16'h3C3D
`define CUBE_LUT_3C15 16'h3C40
`define CUBE_LUT_3C16 16'h3C43
`define CUBE_LUT_3C17 16'h3C47
`define CUBE_LUT_3C18 16'h3C4A
`define CUBE_LUT_3C19 16'h3C4D
`define CUBE_LUT_3C1A 16'h3C50
`define CUBE_LUT_3C1B 16'h3C53
`define CUBE_LUT_3C1C 16'h3C56
`define CUBE_LUT_3C1D 16'h3C59
`define CUBE_LUT_3C1E 16'h3C5D
`define CUBE_LUT_3C1F 16'h3C60
`define CUBE_LUT_3C20 16'h3C63
`define CUBE_LUT_3C21 16'h3C66
`define CUBE_LUT_3C22 16'h3C69
`define CUBE_LUT_3C23 16'h3C6D
`define CUBE_LUT_3C24 16'h3C70
`define CUBE_LUT_3C25 16'h3C73
`define CUBE_LUT_3C26 16'h3C76
`define CUBE_LUT_3C27 16'h3C7A
`define CUBE_LUT_3C28 16'h3C7D
`define CUBE_LUT_3C29 16'h3C80
`define CUBE_LUT_3C2A 16'h3C83
`define CUBE_LUT_3C2B 16'h3C86
`define CUBE_LUT_3C2C 16'h3C8A
`define CUBE_LUT_3C2D 16'h3C8D
`define CUBE_LUT_3C2E 16'h3C90
`define CUBE_LUT_3C2F 16'h3C94
`define CUBE_LUT_3C30 16'h3C97
`define CUBE_LUT_3C31 16'h3C9A
`define CUBE_LUT_3C32 16'h3C9D
`define CUBE_LUT_3C33 16'h3CA1
`define CUBE_LUT_3C34 16'h3CA4
`define CUBE_LUT_3C35 16'h3CA7
`define CUBE_LUT_3C36 16'h3CAB
`define CUBE_LUT_3C37 16'h3CAE
`define CUBE_LUT_3C38 16'h3CB1
`define CUBE_LUT_3C39 16'h3CB5
`define CUBE_LUT_3C3A 16'h3CB8
`define CUBE_LUT_3C3B 16'h3CBB
`define CUBE_LUT_3C3C 16'h3CBF
`define CUBE_LUT_3C3D 16'h3CC2
`define CUBE_LUT_3C3E 16'h3CC5
`define CUBE_LUT_3C3F 16'h3CC9
`define CUBE_LUT_3C40 16'h3CCC
`define CUBE_LUT_3C41 16'h3CD0
`define CUBE_LUT_3C42 16'h3CD3
`define CUBE_LUT_3C43 16'h3CD6
`define CUBE_LUT_3C44 16'h3CDA
`define CUBE_LUT_3C45 16'h3CDD
`define CUBE_LUT_3C46 16'h3CE1
`define CUBE_LUT_3C47 16'h3CE4
`define CUBE_LUT_3C48 16'h3CE8
`define CUBE_LUT_3C49 16'h3CEB
`define CUBE_LUT_3C4A 16'h3CEE
`define CUBE_LUT_3C4B 16'h3CF2
`define CUBE_LUT_3C4C 16'h3CF5
`define CUBE_LUT_3C4D 16'h3CF9
`define CUBE_LUT_3C4E 16'h3CFC
`define CUBE_LUT_3C4F 16'h3D00
`define CUBE_LUT_3C50 16'h3D03
`define CUBE_LUT_3C51 16'h3D07
`define CUBE_LUT_3C52 16'h3D0A
`define CUBE_LUT_3C53 16'h3D0E
`define CUBE_LUT_3C54 16'h3D11
`define CUBE_LUT_3C55 16'h3D15
`define CUBE_LUT_3C56 16'h3D18
`define CUBE_LUT_3C57 16'h3D1C
`define CUBE_LUT_3C58 16'h3D1F
`define CUBE_LUT_3C59 16'h3D23
`define CUBE_LUT_3C5A 16'h3D26
`define CUBE_LUT_3C5B 16'h3D2A
`define CUBE_LUT_3C5C 16'h3D2E
`define CUBE_LUT_3C5D 16'h3D31
`define CUBE_LUT_3C5E 16'h3D35
`define CUBE_LUT_3C5F 16'h3D38
`define CUBE_LUT_3C60 16'h3D3C
`define CUBE_LUT_3C61 16'h3D3F
`define CUBE_LUT_3C62 16'h3D43
`define CUBE_LUT_3C63 16'h3D47
`define CUBE_LUT_3C64 16'h3D4A
`define CUBE_LUT_3C65 16'h3D4E
`define CUBE_LUT_3C66 16'h3D51
`define CUBE_LUT_3C67 16'h3D55
`define CUBE_LUT_3C68 16'h3D59
`define CUBE_LUT_3C69 16'h3D5C
`define CUBE_LUT_3C6A 16'h3D60
`define CUBE_LUT_3C6B 16'h3D64
`define CUBE_LUT_3C6C 16'h3D67
`define CUBE_LUT_3C6D 16'h3D6B
`define CUBE_LUT_3C6E 16'h3D6F
`define CUBE_LUT_3C6F 16'h3D72
`define CUBE_LUT_3C70 16'h3D76
`define CUBE_LUT_3C71 16'h3D7A
`define CUBE_LUT_3C72 16'h3D7D
`define CUBE_LUT_3C73 16'h3D81
`define CUBE_LUT_3C74 16'h3D85
`define CUBE_LUT_3C75 16'h3D89
`define CUBE_LUT_3C76 16'h3D8C
`define CUBE_LUT_3C77 16'h3D90
`define CUBE_LUT_3C78 16'h3D94
`define CUBE_LUT_3C79 16'h3D98
`define CUBE_LUT_3C7A 16'h3D9B
`define CUBE_LUT_3C7B 16'h3D9F
`define CUBE_LUT_3C7C 16'h3DA3
`define CUBE_LUT_3C7D 16'h3DA7
`define CUBE_LUT_3C7E 16'h3DAA
`define CUBE_LUT_3C7F 16'h3DAE
`define CUBE_LUT_3C80 16'h3DB2
`define CUBE_LUT_3C81 16'h3DB6
`define CUBE_LUT_3C82 16'h3DBA
`define CUBE_LUT_3C83 16'h3DBD
`define CUBE_LUT_3C84 16'h3DC1
`define CUBE_LUT_3C85 16'h3DC5
`define CUBE_LUT_3C86 16'h3DC9
`define CUBE_LUT_3C87 16'h3DCD
`define CUBE_LUT_3C88 16'h3DD1
`define CUBE_LUT_3C89 16'h3DD4
`define CUBE_LUT_3C8A 16'h3DD8
`define CUBE_LUT_3C8B 16'h3DDC
`define CUBE_LUT_3C8C 16'h3DE0
`define CUBE_LUT_3C8D 16'h3DE4
`define CUBE_LUT_3C8E 16'h3DE8
`define CUBE_LUT_3C8F 16'h3DEC
`define CUBE_LUT_3C90 16'h3DF0
`define CUBE_LUT_3C91 16'h3DF4
`define CUBE_LUT_3C92 16'h3DF7
`define CUBE_LUT_3C93 16'h3DFB
`define CUBE_LUT_3C94 16'h3DFF
`define CUBE_LUT_3C95 16'h3E03
`define CUBE_LUT_3C96 16'h3E07
`define CUBE_LUT_3C97 16'h3E0B
`define CUBE_LUT_3C98 16'h3E0F
`define CUBE_LUT_3C99 16'h3E13
`define CUBE_LUT_3C9A 16'h3E17
`define CUBE_LUT_3C9B 16'h3E1B
`define CUBE_LUT_3C9C 16'h3E1F
`define CUBE_LUT_3C9D 16'h3E23
`define CUBE_LUT_3C9E 16'h3E27
`define CUBE_LUT_3C9F 16'h3E2B
`define CUBE_LUT_3CA0 16'h3E2F
`define CUBE_LUT_3CA1 16'h3E33
`define CUBE_LUT_3CA2 16'h3E37
`define CUBE_LUT_3CA3 16'h3E3B
`define CUBE_LUT_3CA4 16'h3E3F
`define CUBE_LUT_3CA5 16'h3E43
`define CUBE_LUT_3CA6 16'h3E47
`define CUBE_LUT_3CA7 16'h3E4B
`define CUBE_LUT_3CA8 16'h3E4F
`define CUBE_LUT_3CA9 16'h3E53
`define CUBE_LUT_3CAA 16'h3E57
`define CUBE_LUT_3CAB 16'h3E5B
`define CUBE_LUT_3CAC 16'h3E60
`define CUBE_LUT_3CAD 16'h3E64
`define CUBE_LUT_3CAE 16'h3E68
`define CUBE_LUT_3CAF 16'h3E6C
`define CUBE_LUT_3CB0 16'h3E70
`define CUBE_LUT_3CB1 16'h3E74
`define CUBE_LUT_3CB2 16'h3E78
`define CUBE_LUT_3CB3 16'h3E7C
`define CUBE_LUT_3CB4 16'h3E80
`define CUBE_LUT_3CB5 16'h3E85
`define CUBE_LUT_3CB6 16'h3E89
`define CUBE_LUT_3CB7 16'h3E8D
`define CUBE_LUT_3CB8 16'h3E91
`define CUBE_LUT_3CB9 16'h3E95
`define CUBE_LUT_3CBA 16'h3E99
`define CUBE_LUT_3CBB 16'h3E9E
`define CUBE_LUT_3CBC 16'h3EA2
`define CUBE_LUT_3CBD 16'h3EA6
`define CUBE_LUT_3CBE 16'h3EAA
`define CUBE_LUT_3CBF 16'h3EAF
`define CUBE_LUT_3CC0 16'h3EB3
`define CUBE_LUT_3CC1 16'h3EB7
`define CUBE_LUT_3CC2 16'h3EBB
`define CUBE_LUT_3CC3 16'h3EBF
`define CUBE_LUT_3CC4 16'h3EC4
`define CUBE_LUT_3CC5 16'h3EC8
`define CUBE_LUT_3CC6 16'h3ECC
`define CUBE_LUT_3CC7 16'h3ED1
`define CUBE_LUT_3CC8 16'h3ED5
`define CUBE_LUT_3CC9 16'h3ED9
`define CUBE_LUT_3CCA 16'h3EDD
`define CUBE_LUT_3CCB 16'h3EE2
`define CUBE_LUT_3CCC 16'h3EE6
`define CUBE_LUT_3CCD 16'h3EEA
`define CUBE_LUT_3CCE 16'h3EEF
`define CUBE_LUT_3CCF 16'h3EF3
`define CUBE_LUT_3CD0 16'h3EF7
`define CUBE_LUT_3CD1 16'h3EFC
`define CUBE_LUT_3CD2 16'h3F00
`define CUBE_LUT_3CD3 16'h3F04
`define CUBE_LUT_3CD4 16'h3F09
`define CUBE_LUT_3CD5 16'h3F0D
`define CUBE_LUT_3CD6 16'h3F12
`define CUBE_LUT_3CD7 16'h3F16
`define CUBE_LUT_3CD8 16'h3F1A
`define CUBE_LUT_3CD9 16'h3F1F
`define CUBE_LUT_3CDA 16'h3F23
`define CUBE_LUT_3CDB 16'h3F28
`define CUBE_LUT_3CDC 16'h3F2C
`define CUBE_LUT_3CDD 16'h3F30
`define CUBE_LUT_3CDE 16'h3F35
`define CUBE_LUT_3CDF 16'h3F39
`define CUBE_LUT_3CE0 16'h3F3E
`define CUBE_LUT_3CE1 16'h3F42
`define CUBE_LUT_3CE2 16'h3F47
`define CUBE_LUT_3CE3 16'h3F4B
`define CUBE_LUT_3CE4 16'h3F50
`define CUBE_LUT_3CE5 16'h3F54
`define CUBE_LUT_3CE6 16'h3F59
`define CUBE_LUT_3CE7 16'h3F5D
`define CUBE_LUT_3CE8 16'h3F62
`define CUBE_LUT_3CE9 16'h3F66
`define CUBE_LUT_3CEA 16'h3F6B
`define CUBE_LUT_3CEB 16'h3F6F
`define CUBE_LUT_3CEC 16'h3F74
`define CUBE_LUT_3CED 16'h3F78
`define CUBE_LUT_3CEE 16'h3F7D
`define CUBE_LUT_3CEF 16'h3F81
`define CUBE_LUT_3CF0 16'h3F86
`define CUBE_LUT_3CF1 16'h3F8B
`define CUBE_LUT_3CF2 16'h3F8F
`define CUBE_LUT_3CF3 16'h3F94
`define CUBE_LUT_3CF4 16'h3F98
`define CUBE_LUT_3CF5 16'h3F9D
`define CUBE_LUT_3CF6 16'h3FA1
`define CUBE_LUT_3CF7 16'h3FA6
`define CUBE_LUT_3CF8 16'h3FAB
`define CUBE_LUT_3CF9 16'h3FAF
`define CUBE_LUT_3CFA 16'h3FB4
`define CUBE_LUT_3CFB 16'h3FB9
`define CUBE_LUT_3CFC 16'h3FBD
`define CUBE_LUT_3CFD 16'h3FC2
`define CUBE_LUT_3CFE 16'h3FC7
`define CUBE_LUT_3CFF 16'h3FCB
`define CUBE_LUT_3D00 16'h3FD0
`define CUBE_LUT_3D01 16'h3FD5
`define CUBE_LUT_3D02 16'h3FD9
`define CUBE_LUT_3D03 16'h3FDE
`define CUBE_LUT_3D04 16'h3FE3
`define CUBE_LUT_3D05 16'h3FE8
`define CUBE_LUT_3D06 16'h3FEC
`define CUBE_LUT_3D07 16'h3FF1
`define CUBE_LUT_3D08 16'h3FF6
`define CUBE_LUT_3D09 16'h3FFA
`define CUBE_LUT_3D0A 16'h3FFF
`define CUBE_LUT_3D0B 16'h4002
`define CUBE_LUT_3D0C 16'h4004
`define CUBE_LUT_3D0D 16'h4007
`define CUBE_LUT_3D0E 16'h4009
`define CUBE_LUT_3D0F 16'h400C
`define CUBE_LUT_3D10 16'h400E
`define CUBE_LUT_3D11 16'h4010
`define CUBE_LUT_3D12 16'h4013
`define CUBE_LUT_3D13 16'h4015
`define CUBE_LUT_3D14 16'h4018
`define CUBE_LUT_3D15 16'h401A
`define CUBE_LUT_3D16 16'h401C
`define CUBE_LUT_3D17 16'h401F
`define CUBE_LUT_3D18 16'h4021
`define CUBE_LUT_3D19 16'h4024
`define CUBE_LUT_3D1A 16'h4026
`define CUBE_LUT_3D1B 16'h4029
`define CUBE_LUT_3D1C 16'h402B
`define CUBE_LUT_3D1D 16'h402E
`define CUBE_LUT_3D1E 16'h4030
`define CUBE_LUT_3D1F 16'h4032
`define CUBE_LUT_3D20 16'h4035
`define CUBE_LUT_3D21 16'h4037
`define CUBE_LUT_3D22 16'h403A
`define CUBE_LUT_3D23 16'h403C
`define CUBE_LUT_3D24 16'h403F
`define CUBE_LUT_3D25 16'h4041
`define CUBE_LUT_3D26 16'h4044
`define CUBE_LUT_3D27 16'h4046
`define CUBE_LUT_3D28 16'h4049
`define CUBE_LUT_3D29 16'h404B
`define CUBE_LUT_3D2A 16'h404E
`define CUBE_LUT_3D2B 16'h4050
`define CUBE_LUT_3D2C 16'h4053
`define CUBE_LUT_3D2D 16'h4055
`define CUBE_LUT_3D2E 16'h4058
`define CUBE_LUT_3D2F 16'h405A
`define CUBE_LUT_3D30 16'h405D
`define CUBE_LUT_3D31 16'h405F
`define CUBE_LUT_3D32 16'h4062
`define CUBE_LUT_3D33 16'h4064
`define CUBE_LUT_3D34 16'h4067
`define CUBE_LUT_3D35 16'h4069
`define CUBE_LUT_3D36 16'h406C
`define CUBE_LUT_3D37 16'h406F
`define CUBE_LUT_3D38 16'h4071
`define CUBE_LUT_3D39 16'h4074
`define CUBE_LUT_3D3A 16'h4076
`define CUBE_LUT_3D3B 16'h4079
`define CUBE_LUT_3D3C 16'h407B
`define CUBE_LUT_3D3D 16'h407E
`define CUBE_LUT_3D3E 16'h4080
`define CUBE_LUT_3D3F 16'h4083
`define CUBE_LUT_3D40 16'h4086
`define CUBE_LUT_3D41 16'h4088
`define CUBE_LUT_3D42 16'h408B
`define CUBE_LUT_3D43 16'h408D
`define CUBE_LUT_3D44 16'h4090
`define CUBE_LUT_3D45 16'h4093
`define CUBE_LUT_3D46 16'h4095
`define CUBE_LUT_3D47 16'h4098
`define CUBE_LUT_3D48 16'h409A
`define CUBE_LUT_3D49 16'h409D
`define CUBE_LUT_3D4A 16'h40A0
`define CUBE_LUT_3D4B 16'h40A2
`define CUBE_LUT_3D4C 16'h40A5
`define CUBE_LUT_3D4D 16'h40A8
`define CUBE_LUT_3D4E 16'h40AA
`define CUBE_LUT_3D4F 16'h40AD
`define CUBE_LUT_3D50 16'h40AF
`define CUBE_LUT_3D51 16'h40B2
`define CUBE_LUT_3D52 16'h40B5
`define CUBE_LUT_3D53 16'h40B7
`define CUBE_LUT_3D54 16'h40BA
`define CUBE_LUT_3D55 16'h40BD
`define CUBE_LUT_3D56 16'h40BF
`define CUBE_LUT_3D57 16'h40C2
`define CUBE_LUT_3D58 16'h40C5
`define CUBE_LUT_3D59 16'h40C7
`define CUBE_LUT_3D5A 16'h40CA
`define CUBE_LUT_3D5B 16'h40CD
`define CUBE_LUT_3D5C 16'h40CF
`define CUBE_LUT_3D5D 16'h40D2
`define CUBE_LUT_3D5E 16'h40D5
`define CUBE_LUT_3D5F 16'h40D8
`define CUBE_LUT_3D60 16'h40DA
`define CUBE_LUT_3D61 16'h40DD
`define CUBE_LUT_3D62 16'h40E0
`define CUBE_LUT_3D63 16'h40E2
`define CUBE_LUT_3D64 16'h40E5
`define CUBE_LUT_3D65 16'h40E8
`define CUBE_LUT_3D66 16'h40EB
`define CUBE_LUT_3D67 16'h40ED
`define CUBE_LUT_3D68 16'h40F0
`define CUBE_LUT_3D69 16'h40F3
`define CUBE_LUT_3D6A 16'h40F6
`define CUBE_LUT_3D6B 16'h40F8
`define CUBE_LUT_3D6C 16'h40FB
`define CUBE_LUT_3D6D 16'h40FE
`define CUBE_LUT_3D6E 16'h4101
`define CUBE_LUT_3D6F 16'h4103
`define CUBE_LUT_3D70 16'h4106
`define CUBE_LUT_3D71 16'h4109
`define CUBE_LUT_3D72 16'h410C
`define CUBE_LUT_3D73 16'h410E
`define CUBE_LUT_3D74 16'h4111
`define CUBE_LUT_3D75 16'h4114
`define CUBE_LUT_3D76 16'h4117
`define CUBE_LUT_3D77 16'h411A
`define CUBE_LUT_3D78 16'h411C
`define CUBE_LUT_3D79 16'h411F
`define CUBE_LUT_3D7A 16'h4122
`define CUBE_LUT_3D7B 16'h4125
`define CUBE_LUT_3D7C 16'h4128
`define CUBE_LUT_3D7D 16'h412B
`define CUBE_LUT_3D7E 16'h412D
`define CUBE_LUT_3D7F 16'h4130
`define CUBE_LUT_3D80 16'h4133
`define CUBE_LUT_3D81 16'h4136
`define CUBE_LUT_3D82 16'h4139
`define CUBE_LUT_3D83 16'h413C
`define CUBE_LUT_3D84 16'h413E
`define CUBE_LUT_3D85 16'h4141
`define CUBE_LUT_3D86 16'h4144
`define CUBE_LUT_3D87 16'h4147
`define CUBE_LUT_3D88 16'h414A
`define CUBE_LUT_3D89 16'h414D
`define CUBE_LUT_3D8A 16'h4150
`define CUBE_LUT_3D8B 16'h4152
`define CUBE_LUT_3D8C 16'h4155
`define CUBE_LUT_3D8D 16'h4158
`define CUBE_LUT_3D8E 16'h415B
`define CUBE_LUT_3D8F 16'h415E
`define CUBE_LUT_3D90 16'h4161
`define CUBE_LUT_3D91 16'h4164
`define CUBE_LUT_3D92 16'h4167
`define CUBE_LUT_3D93 16'h416A
`define CUBE_LUT_3D94 16'h416D
`define CUBE_LUT_3D95 16'h416F
`define CUBE_LUT_3D96 16'h4172
`define CUBE_LUT_3D97 16'h4175
`define CUBE_LUT_3D98 16'h4178
`define CUBE_LUT_3D99 16'h417B
`define CUBE_LUT_3D9A 16'h417E
`define CUBE_LUT_3D9B 16'h4181
`define CUBE_LUT_3D9C 16'h4184
`define CUBE_LUT_3D9D 16'h4187
`define CUBE_LUT_3D9E 16'h418A
`define CUBE_LUT_3D9F 16'h418D
`define CUBE_LUT_3DA0 16'h4190
`define CUBE_LUT_3DA1 16'h4193
`define CUBE_LUT_3DA2 16'h4196
`define CUBE_LUT_3DA3 16'h4199
`define CUBE_LUT_3DA4 16'h419C
`define CUBE_LUT_3DA5 16'h419F
`define CUBE_LUT_3DA6 16'h41A2
`define CUBE_LUT_3DA7 16'h41A5
`define CUBE_LUT_3DA8 16'h41A8
`define CUBE_LUT_3DA9 16'h41AB
`define CUBE_LUT_3DAA 16'h41AE
`define CUBE_LUT_3DAB 16'h41B1
`define CUBE_LUT_3DAC 16'h41B4
`define CUBE_LUT_3DAD 16'h41B7
`define CUBE_LUT_3DAE 16'h41BA
`define CUBE_LUT_3DAF 16'h41BD
`define CUBE_LUT_3DB0 16'h41C0
`define CUBE_LUT_3DB1 16'h41C3
`define CUBE_LUT_3DB2 16'h41C6
`define CUBE_LUT_3DB3 16'h41C9
`define CUBE_LUT_3DB4 16'h41CC
`define CUBE_LUT_3DB5 16'h41CF
`define CUBE_LUT_3DB6 16'h41D2
`define CUBE_LUT_3DB7 16'h41D5
`define CUBE_LUT_3DB8 16'h41D8
`define CUBE_LUT_3DB9 16'h41DB
`define CUBE_LUT_3DBA 16'h41DE
`define CUBE_LUT_3DBB 16'h41E1
`define CUBE_LUT_3DBC 16'h41E5
`define CUBE_LUT_3DBD 16'h41E8
`define CUBE_LUT_3DBE 16'h41EB
`define CUBE_LUT_3DBF 16'h41EE
`define CUBE_LUT_3DC0 16'h41F1
`define CUBE_LUT_3DC1 16'h41F4
`define CUBE_LUT_3DC2 16'h41F7
`define CUBE_LUT_3DC3 16'h41FA
`define CUBE_LUT_3DC4 16'h41FD
`define CUBE_LUT_3DC5 16'h4200
`define CUBE_LUT_3DC6 16'h4204
`define CUBE_LUT_3DC7 16'h4207
`define CUBE_LUT_3DC8 16'h420A
`define CUBE_LUT_3DC9 16'h420D
`define CUBE_LUT_3DCA 16'h4210
`define CUBE_LUT_3DCB 16'h4213
`define CUBE_LUT_3DCC 16'h4216
`define CUBE_LUT_3DCD 16'h421A
`define CUBE_LUT_3DCE 16'h421D
`define CUBE_LUT_3DCF 16'h4220
`define CUBE_LUT_3DD0 16'h4223
`define CUBE_LUT_3DD1 16'h4226
`define CUBE_LUT_3DD2 16'h4229
`define CUBE_LUT_3DD3 16'h422D
`define CUBE_LUT_3DD4 16'h4230
`define CUBE_LUT_3DD5 16'h4233
`define CUBE_LUT_3DD6 16'h4236
`define CUBE_LUT_3DD7 16'h4239
`define CUBE_LUT_3DD8 16'h423C
`define CUBE_LUT_3DD9 16'h4240
`define CUBE_LUT_3DDA 16'h4243
`define CUBE_LUT_3DDB 16'h4246
`define CUBE_LUT_3DDC 16'h4249
`define CUBE_LUT_3DDD 16'h424D
`define CUBE_LUT_3DDE 16'h4250
`define CUBE_LUT_3DDF 16'h4253
`define CUBE_LUT_3DE0 16'h4256
`define CUBE_LUT_3DE1 16'h4259
`define CUBE_LUT_3DE2 16'h425D
`define CUBE_LUT_3DE3 16'h4260
`define CUBE_LUT_3DE4 16'h4263
`define CUBE_LUT_3DE5 16'h4266
`define CUBE_LUT_3DE6 16'h426A
`define CUBE_LUT_3DE7 16'h426D
`define CUBE_LUT_3DE8 16'h4270
`define CUBE_LUT_3DE9 16'h4274
`define CUBE_LUT_3DEA 16'h4277
`define CUBE_LUT_3DEB 16'h427A
`define CUBE_LUT_3DEC 16'h427D
`define CUBE_LUT_3DED 16'h4281
`define CUBE_LUT_3DEE 16'h4284
`define CUBE_LUT_3DEF 16'h4287
`define CUBE_LUT_3DF0 16'h428B
`define CUBE_LUT_3DF1 16'h428E
`define CUBE_LUT_3DF2 16'h4291
`define CUBE_LUT_3DF3 16'h4294
`define CUBE_LUT_3DF4 16'h4298
`define CUBE_LUT_3DF5 16'h429B
`define CUBE_LUT_3DF6 16'h429E
`define CUBE_LUT_3DF7 16'h42A2
`define CUBE_LUT_3DF8 16'h42A5
`define CUBE_LUT_3DF9 16'h42A8
`define CUBE_LUT_3DFA 16'h42AC
`define CUBE_LUT_3DFB 16'h42AF
`define CUBE_LUT_3DFC 16'h42B3
`define CUBE_LUT_3DFD 16'h42B6
`define CUBE_LUT_3DFE 16'h42B9
`define CUBE_LUT_3DFF 16'h42BD
`define CUBE_LUT_3E00 16'h42C0
`define CUBE_LUT_3E01 16'h42C3
`define CUBE_LUT_3E02 16'h42C7
`define CUBE_LUT_3E03 16'h42CA
`define CUBE_LUT_3E04 16'h42CE
`define CUBE_LUT_3E05 16'h42D1
`define CUBE_LUT_3E06 16'h42D4
`define CUBE_LUT_3E07 16'h42D8
`define CUBE_LUT_3E08 16'h42DB
`define CUBE_LUT_3E09 16'h42DF
`define CUBE_LUT_3E0A 16'h42E2
`define CUBE_LUT_3E0B 16'h42E5
`define CUBE_LUT_3E0C 16'h42E9
`define CUBE_LUT_3E0D 16'h42EC
`define CUBE_LUT_3E0E 16'h42F0
`define CUBE_LUT_3E0F 16'h42F3
`define CUBE_LUT_3E10 16'h42F7
`define CUBE_LUT_3E11 16'h42FA
`define CUBE_LUT_3E12 16'h42FD
`define CUBE_LUT_3E13 16'h4301
`define CUBE_LUT_3E14 16'h4304
`define CUBE_LUT_3E15 16'h4308
`define CUBE_LUT_3E16 16'h430B
`define CUBE_LUT_3E17 16'h430F
`define CUBE_LUT_3E18 16'h4312
`define CUBE_LUT_3E19 16'h4316
`define CUBE_LUT_3E1A 16'h4319
`define CUBE_LUT_3E1B 16'h431D
`define CUBE_LUT_3E1C 16'h4320
`define CUBE_LUT_3E1D 16'h4324
`define CUBE_LUT_3E1E 16'h4327
`define CUBE_LUT_3E1F 16'h432B
`define CUBE_LUT_3E20 16'h432E
`define CUBE_LUT_3E21 16'h4332
`define CUBE_LUT_3E22 16'h4335
`define CUBE_LUT_3E23 16'h4339
`define CUBE_LUT_3E24 16'h433C
`define CUBE_LUT_3E25 16'h4340
`define CUBE_LUT_3E26 16'h4343
`define CUBE_LUT_3E27 16'h4347
`define CUBE_LUT_3E28 16'h434B
`define CUBE_LUT_3E29 16'h434E
`define CUBE_LUT_3E2A 16'h4352
`define CUBE_LUT_3E2B 16'h4355
`define CUBE_LUT_3E2C 16'h4359
`define CUBE_LUT_3E2D 16'h435C
`define CUBE_LUT_3E2E 16'h4360
`define CUBE_LUT_3E2F 16'h4364
`define CUBE_LUT_3E30 16'h4367
`define CUBE_LUT_3E31 16'h436B
`define CUBE_LUT_3E32 16'h436E
`define CUBE_LUT_3E33 16'h4372
`define CUBE_LUT_3E34 16'h4376
`define CUBE_LUT_3E35 16'h4379
`define CUBE_LUT_3E36 16'h437D
`define CUBE_LUT_3E37 16'h4380
`define CUBE_LUT_3E38 16'h4384
`define CUBE_LUT_3E39 16'h4388
`define CUBE_LUT_3E3A 16'h438B
`define CUBE_LUT_3E3B 16'h438F
`define CUBE_LUT_3E3C 16'h4393
`define CUBE_LUT_3E3D 16'h4396
`define CUBE_LUT_3E3E 16'h439A
`define CUBE_LUT_3E3F 16'h439D
`define CUBE_LUT_3E40 16'h43A1
`define CUBE_LUT_3E41 16'h43A5
`define CUBE_LUT_3E42 16'h43A8
`define CUBE_LUT_3E43 16'h43AC
`define CUBE_LUT_3E44 16'h43B0
`define CUBE_LUT_3E45 16'h43B3
`define CUBE_LUT_3E46 16'h43B7
`define CUBE_LUT_3E47 16'h43BB
`define CUBE_LUT_3E48 16'h43BF
`define CUBE_LUT_3E49 16'h43C2
`define CUBE_LUT_3E4A 16'h43C6
`define CUBE_LUT_3E4B 16'h43CA
`define CUBE_LUT_3E4C 16'h43CD
`define CUBE_LUT_3E4D 16'h43D1
`define CUBE_LUT_3E4E 16'h43D5
`define CUBE_LUT_3E4F 16'h43D9
`define CUBE_LUT_3E50 16'h43DC
`define CUBE_LUT_3E51 16'h43E0
`define CUBE_LUT_3E52 16'h43E4
`define CUBE_LUT_3E53 16'h43E8
`define CUBE_LUT_3E54 16'h43EB
`define CUBE_LUT_3E55 16'h43EF
`define CUBE_LUT_3E56 16'h43F3
`define CUBE_LUT_3E57 16'h43F7
`define CUBE_LUT_3E58 16'h43FA
`define CUBE_LUT_3E59 16'h43FE
`define CUBE_LUT_3E5A 16'h4401
`define CUBE_LUT_3E5B 16'h4403
`define CUBE_LUT_3E5C 16'h4405
`define CUBE_LUT_3E5D 16'h4407
`define CUBE_LUT_3E5E 16'h4409
`define CUBE_LUT_3E5F 16'h440A
`define CUBE_LUT_3E60 16'h440C
`define CUBE_LUT_3E61 16'h440E
`define CUBE_LUT_3E62 16'h4410
`define CUBE_LUT_3E63 16'h4412
`define CUBE_LUT_3E64 16'h4414
`define CUBE_LUT_3E65 16'h4416
`define CUBE_LUT_3E66 16'h4418
`define CUBE_LUT_3E67 16'h441A
`define CUBE_LUT_3E68 16'h441C
`define CUBE_LUT_3E69 16'h441E
`define CUBE_LUT_3E6A 16'h4420
`define CUBE_LUT_3E6B 16'h4421
`define CUBE_LUT_3E6C 16'h4423
`define CUBE_LUT_3E6D 16'h4425
`define CUBE_LUT_3E6E 16'h4427
`define CUBE_LUT_3E6F 16'h4429
`define CUBE_LUT_3E70 16'h442B
`define CUBE_LUT_3E71 16'h442D
`define CUBE_LUT_3E72 16'h442F
`define CUBE_LUT_3E73 16'h4431
`define CUBE_LUT_3E74 16'h4433
`define CUBE_LUT_3E75 16'h4435
`define CUBE_LUT_3E76 16'h4437
`define CUBE_LUT_3E77 16'h4439
`define CUBE_LUT_3E78 16'h443B
`define CUBE_LUT_3E79 16'h443D
`define CUBE_LUT_3E7A 16'h443F
`define CUBE_LUT_3E7B 16'h4441
`define CUBE_LUT_3E7C 16'h4443
`define CUBE_LUT_3E7D 16'h4445
`define CUBE_LUT_3E7E 16'h4447
`define CUBE_LUT_3E7F 16'h4449
`define CUBE_LUT_3E80 16'h444A
`define CUBE_LUT_3E81 16'h444C
`define CUBE_LUT_3E82 16'h444E
`define CUBE_LUT_3E83 16'h4450
`define CUBE_LUT_3E84 16'h4452
`define CUBE_LUT_3E85 16'h4454
`define CUBE_LUT_3E86 16'h4456
`define CUBE_LUT_3E87 16'h4458
`define CUBE_LUT_3E88 16'h445A
`define CUBE_LUT_3E89 16'h445C
`define CUBE_LUT_3E8A 16'h445E
`define CUBE_LUT_3E8B 16'h4460
`define CUBE_LUT_3E8C 16'h4462
`define CUBE_LUT_3E8D 16'h4464
`define CUBE_LUT_3E8E 16'h4466
`define CUBE_LUT_3E8F 16'h4468
`define CUBE_LUT_3E90 16'h446A
`define CUBE_LUT_3E91 16'h446D
`define CUBE_LUT_3E92 16'h446F
`define CUBE_LUT_3E93 16'h4471
`define CUBE_LUT_3E94 16'h4473
`define CUBE_LUT_3E95 16'h4475
`define CUBE_LUT_3E96 16'h4477
`define CUBE_LUT_3E97 16'h4479
`define CUBE_LUT_3E98 16'h447B
`define CUBE_LUT_3E99 16'h447D
`define CUBE_LUT_3E9A 16'h447F
`define CUBE_LUT_3E9B 16'h4481
`define CUBE_LUT_3E9C 16'h4483
`define CUBE_LUT_3E9D 16'h4485
`define CUBE_LUT_3E9E 16'h4487
`define CUBE_LUT_3E9F 16'h4489
`define CUBE_LUT_3EA0 16'h448B
`define CUBE_LUT_3EA1 16'h448D
`define CUBE_LUT_3EA2 16'h448F
`define CUBE_LUT_3EA3 16'h4491
`define CUBE_LUT_3EA4 16'h4493
`define CUBE_LUT_3EA5 16'h4495
`define CUBE_LUT_3EA6 16'h4497
`define CUBE_LUT_3EA7 16'h449A
`define CUBE_LUT_3EA8 16'h449C
`define CUBE_LUT_3EA9 16'h449E
`define CUBE_LUT_3EAA 16'h44A0
`define CUBE_LUT_3EAB 16'h44A2
`define CUBE_LUT_3EAC 16'h44A4
`define CUBE_LUT_3EAD 16'h44A6
`define CUBE_LUT_3EAE 16'h44A8
`define CUBE_LUT_3EAF 16'h44AA
`define CUBE_LUT_3EB0 16'h44AC
`define CUBE_LUT_3EB1 16'h44AE
`define CUBE_LUT_3EB2 16'h44B1
`define CUBE_LUT_3EB3 16'h44B3
`define CUBE_LUT_3EB4 16'h44B5
`define CUBE_LUT_3EB5 16'h44B7
`define CUBE_LUT_3EB6 16'h44B9
`define CUBE_LUT_3EB7 16'h44BB
`define CUBE_LUT_3EB8 16'h44BD
`define CUBE_LUT_3EB9 16'h44BF
`define CUBE_LUT_3EBA 16'h44C1
`define CUBE_LUT_3EBB 16'h44C4
`define CUBE_LUT_3EBC 16'h44C6
`define CUBE_LUT_3EBD 16'h44C8
`define CUBE_LUT_3EBE 16'h44CA
`define CUBE_LUT_3EBF 16'h44CC
`define CUBE_LUT_3EC0 16'h44CE
`define CUBE_LUT_3EC1 16'h44D0
`define CUBE_LUT_3EC2 16'h44D2
`define CUBE_LUT_3EC3 16'h44D5
`define CUBE_LUT_3EC4 16'h44D7
`define CUBE_LUT_3EC5 16'h44D9
`define CUBE_LUT_3EC6 16'h44DB
`define CUBE_LUT_3EC7 16'h44DD
`define CUBE_LUT_3EC8 16'h44DF
`define CUBE_LUT_3EC9 16'h44E2
`define CUBE_LUT_3ECA 16'h44E4
`define CUBE_LUT_3ECB 16'h44E6
`define CUBE_LUT_3ECC 16'h44E8
`define CUBE_LUT_3ECD 16'h44EA
`define CUBE_LUT_3ECE 16'h44EC
`define CUBE_LUT_3ECF 16'h44EF
`define CUBE_LUT_3ED0 16'h44F1
`define CUBE_LUT_3ED1 16'h44F3
`define CUBE_LUT_3ED2 16'h44F5
`define CUBE_LUT_3ED3 16'h44F7
`define CUBE_LUT_3ED4 16'h44F9
`define CUBE_LUT_3ED5 16'h44FC
`define CUBE_LUT_3ED6 16'h44FE
`define CUBE_LUT_3ED7 16'h4500
`define CUBE_LUT_3ED8 16'h4502
`define CUBE_LUT_3ED9 16'h4504
`define CUBE_LUT_3EDA 16'h4507
`define CUBE_LUT_3EDB 16'h4509
`define CUBE_LUT_3EDC 16'h450B
`define CUBE_LUT_3EDD 16'h450D
`define CUBE_LUT_3EDE 16'h450F
`define CUBE_LUT_3EDF 16'h4512
`define CUBE_LUT_3EE0 16'h4514
`define CUBE_LUT_3EE1 16'h4516
`define CUBE_LUT_3EE2 16'h4518
`define CUBE_LUT_3EE3 16'h451A
`define CUBE_LUT_3EE4 16'h451D
`define CUBE_LUT_3EE5 16'h451F
`define CUBE_LUT_3EE6 16'h4521
`define CUBE_LUT_3EE7 16'h4523
`define CUBE_LUT_3EE8 16'h4526
`define CUBE_LUT_3EE9 16'h4528
`define CUBE_LUT_3EEA 16'h452A
`define CUBE_LUT_3EEB 16'h452C
`define CUBE_LUT_3EEC 16'h452F
`define CUBE_LUT_3EED 16'h4531
`define CUBE_LUT_3EEE 16'h4533
`define CUBE_LUT_3EEF 16'h4535
`define CUBE_LUT_3EF0 16'h4538
`define CUBE_LUT_3EF1 16'h453A
`define CUBE_LUT_3EF2 16'h453C
`define CUBE_LUT_3EF3 16'h453E
`define CUBE_LUT_3EF4 16'h4541
`define CUBE_LUT_3EF5 16'h4543
`define CUBE_LUT_3EF6 16'h4545
`define CUBE_LUT_3EF7 16'h4547
`define CUBE_LUT_3EF8 16'h454A
`define CUBE_LUT_3EF9 16'h454C
`define CUBE_LUT_3EFA 16'h454E
`define CUBE_LUT_3EFB 16'h4551
`define CUBE_LUT_3EFC 16'h4553
`define CUBE_LUT_3EFD 16'h4555
`define CUBE_LUT_3EFE 16'h4557
`define CUBE_LUT_3EFF 16'h455A
`define CUBE_LUT_3F00 16'h455C
`define CUBE_LUT_3F01 16'h455E
`define CUBE_LUT_3F02 16'h4561
`define CUBE_LUT_3F03 16'h4563
`define CUBE_LUT_3F04 16'h4565
`define CUBE_LUT_3F05 16'h4568
`define CUBE_LUT_3F06 16'h456A
`define CUBE_LUT_3F07 16'h456C
`define CUBE_LUT_3F08 16'h456E
`define CUBE_LUT_3F09 16'h4571
`define CUBE_LUT_3F0A 16'h4573
`define CUBE_LUT_3F0B 16'h4575
`define CUBE_LUT_3F0C 16'h4578
`define CUBE_LUT_3F0D 16'h457A
`define CUBE_LUT_3F0E 16'h457C
`define CUBE_LUT_3F0F 16'h457F
`define CUBE_LUT_3F10 16'h4581
`define CUBE_LUT_3F11 16'h4583
`define CUBE_LUT_3F12 16'h4586
`define CUBE_LUT_3F13 16'h4588
`define CUBE_LUT_3F14 16'h458A
`define CUBE_LUT_3F15 16'h458D
`define CUBE_LUT_3F16 16'h458F
`define CUBE_LUT_3F17 16'h4592
`define CUBE_LUT_3F18 16'h4594
`define CUBE_LUT_3F19 16'h4596
`define CUBE_LUT_3F1A 16'h4599
`define CUBE_LUT_3F1B 16'h459B
`define CUBE_LUT_3F1C 16'h459D
`define CUBE_LUT_3F1D 16'h45A0
`define CUBE_LUT_3F1E 16'h45A2
`define CUBE_LUT_3F1F 16'h45A4
`define CUBE_LUT_3F20 16'h45A7
`define CUBE_LUT_3F21 16'h45A9
`define CUBE_LUT_3F22 16'h45AC
`define CUBE_LUT_3F23 16'h45AE
`define CUBE_LUT_3F24 16'h45B0
`define CUBE_LUT_3F25 16'h45B3
`define CUBE_LUT_3F26 16'h45B5
`define CUBE_LUT_3F27 16'h45B8
`define CUBE_LUT_3F28 16'h45BA
`define CUBE_LUT_3F29 16'h45BC
`define CUBE_LUT_3F2A 16'h45BF
`define CUBE_LUT_3F2B 16'h45C1
`define CUBE_LUT_3F2C 16'h45C4
`define CUBE_LUT_3F2D 16'h45C6
`define CUBE_LUT_3F2E 16'h45C8
`define CUBE_LUT_3F2F 16'h45CB
`define CUBE_LUT_3F30 16'h45CD
`define CUBE_LUT_3F31 16'h45D0
`define CUBE_LUT_3F32 16'h45D2
`define CUBE_LUT_3F33 16'h45D5
`define CUBE_LUT_3F34 16'h45D7
`define CUBE_LUT_3F35 16'h45D9
`define CUBE_LUT_3F36 16'h45DC
`define CUBE_LUT_3F37 16'h45DE
`define CUBE_LUT_3F38 16'h45E1
`define CUBE_LUT_3F39 16'h45E3
`define CUBE_LUT_3F3A 16'h45E6
`define CUBE_LUT_3F3B 16'h45E8
`define CUBE_LUT_3F3C 16'h45EA
`define CUBE_LUT_3F3D 16'h45ED
`define CUBE_LUT_3F3E 16'h45EF
`define CUBE_LUT_3F3F 16'h45F2
`define CUBE_LUT_3F40 16'h45F4
`define CUBE_LUT_3F41 16'h45F7
`define CUBE_LUT_3F42 16'h45F9
`define CUBE_LUT_3F43 16'h45FC
`define CUBE_LUT_3F44 16'h45FE
`define CUBE_LUT_3F45 16'h4601
`define CUBE_LUT_3F46 16'h4603
`define CUBE_LUT_3F47 16'h4606
`define CUBE_LUT_3F48 16'h4608
`define CUBE_LUT_3F49 16'h460B
`define CUBE_LUT_3F4A 16'h460D
`define CUBE_LUT_3F4B 16'h4610
`define CUBE_LUT_3F4C 16'h4612
`define CUBE_LUT_3F4D 16'h4615
`define CUBE_LUT_3F4E 16'h4617
`define CUBE_LUT_3F4F 16'h461A
`define CUBE_LUT_3F50 16'h461C
`define CUBE_LUT_3F51 16'h461F
`define CUBE_LUT_3F52 16'h4621
`define CUBE_LUT_3F53 16'h4624
`define CUBE_LUT_3F54 16'h4626
`define CUBE_LUT_3F55 16'h4629
`define CUBE_LUT_3F56 16'h462B
`define CUBE_LUT_3F57 16'h462E
`define CUBE_LUT_3F58 16'h4630
`define CUBE_LUT_3F59 16'h4633
`define CUBE_LUT_3F5A 16'h4635
`define CUBE_LUT_3F5B 16'h4638
`define CUBE_LUT_3F5C 16'h463A
`define CUBE_LUT_3F5D 16'h463D
`define CUBE_LUT_3F5E 16'h463F
`define CUBE_LUT_3F5F 16'h4642
`define CUBE_LUT_3F60 16'h4645
`define CUBE_LUT_3F61 16'h4647
`define CUBE_LUT_3F62 16'h464A
`define CUBE_LUT_3F63 16'h464C
`define CUBE_LUT_3F64 16'h464F
`define CUBE_LUT_3F65 16'h4651
`define CUBE_LUT_3F66 16'h4654
`define CUBE_LUT_3F67 16'h4656
`define CUBE_LUT_3F68 16'h4659
`define CUBE_LUT_3F69 16'h465C
`define CUBE_LUT_3F6A 16'h465E
`define CUBE_LUT_3F6B 16'h4661
`define CUBE_LUT_3F6C 16'h4663
`define CUBE_LUT_3F6D 16'h4666
`define CUBE_LUT_3F6E 16'h4668
`define CUBE_LUT_3F6F 16'h466B
`define CUBE_LUT_3F70 16'h466E
`define CUBE_LUT_3F71 16'h4670
`define CUBE_LUT_3F72 16'h4673
`define CUBE_LUT_3F73 16'h4675
`define CUBE_LUT_3F74 16'h4678
`define CUBE_LUT_3F75 16'h467B
`define CUBE_LUT_3F76 16'h467D
`define CUBE_LUT_3F77 16'h4680
`define CUBE_LUT_3F78 16'h4682
`define CUBE_LUT_3F79 16'h4685
`define CUBE_LUT_3F7A 16'h4688
`define CUBE_LUT_3F7B 16'h468A
`define CUBE_LUT_3F7C 16'h468D
`define CUBE_LUT_3F7D 16'h4690
`define CUBE_LUT_3F7E 16'h4692
`define CUBE_LUT_3F7F 16'h4695
`define CUBE_LUT_3F80 16'h4698
`define CUBE_LUT_3F81 16'h469A
`define CUBE_LUT_3F82 16'h469D
`define CUBE_LUT_3F83 16'h469F
`define CUBE_LUT_3F84 16'h46A2
`define CUBE_LUT_3F85 16'h46A5
`define CUBE_LUT_3F86 16'h46A7
`define CUBE_LUT_3F87 16'h46AA
`define CUBE_LUT_3F88 16'h46AD
`define CUBE_LUT_3F89 16'h46AF
`define CUBE_LUT_3F8A 16'h46B2
`define CUBE_LUT_3F8B 16'h46B5
`define CUBE_LUT_3F8C 16'h46B7
`define CUBE_LUT_3F8D 16'h46BA
`define CUBE_LUT_3F8E 16'h46BD
`define CUBE_LUT_3F8F 16'h46BF
`define CUBE_LUT_3F90 16'h46C2
`define CUBE_LUT_3F91 16'h46C5
`define CUBE_LUT_3F92 16'h46C7
`define CUBE_LUT_3F93 16'h46CA
`define CUBE_LUT_3F94 16'h46CD
`define CUBE_LUT_3F95 16'h46CF
`define CUBE_LUT_3F96 16'h46D2
`define CUBE_LUT_3F97 16'h46D5
`define CUBE_LUT_3F98 16'h46D8
`define CUBE_LUT_3F99 16'h46DA
`define CUBE_LUT_3F9A 16'h46DD
`define CUBE_LUT_3F9B 16'h46E0
`define CUBE_LUT_3F9C 16'h46E2
`define CUBE_LUT_3F9D 16'h46E5
`define CUBE_LUT_3F9E 16'h46E8
`define CUBE_LUT_3F9F 16'h46EB
`define CUBE_LUT_3FA0 16'h46ED
`define CUBE_LUT_3FA1 16'h46F0
`define CUBE_LUT_3FA2 16'h46F3
`define CUBE_LUT_3FA3 16'h46F5
`define CUBE_LUT_3FA4 16'h46F8
`define CUBE_LUT_3FA5 16'h46FB
`define CUBE_LUT_3FA6 16'h46FE
`define CUBE_LUT_3FA7 16'h4700
`define CUBE_LUT_3FA8 16'h4703
`define CUBE_LUT_3FA9 16'h4706
`define CUBE_LUT_3FAA 16'h4709
`define CUBE_LUT_3FAB 16'h470B
`define CUBE_LUT_3FAC 16'h470E
`define CUBE_LUT_3FAD 16'h4711
`define CUBE_LUT_3FAE 16'h4714
`define CUBE_LUT_3FAF 16'h4716
`define CUBE_LUT_3FB0 16'h4719
`define CUBE_LUT_3FB1 16'h471C
`define CUBE_LUT_3FB2 16'h471F
`define CUBE_LUT_3FB3 16'h4722
`define CUBE_LUT_3FB4 16'h4724
`define CUBE_LUT_3FB5 16'h4727
`define CUBE_LUT_3FB6 16'h472A
`define CUBE_LUT_3FB7 16'h472D
`define CUBE_LUT_3FB8 16'h4730
`define CUBE_LUT_3FB9 16'h4732
`define CUBE_LUT_3FBA 16'h4735
`define CUBE_LUT_3FBB 16'h4738
`define CUBE_LUT_3FBC 16'h473B
`define CUBE_LUT_3FBD 16'h473E
`define CUBE_LUT_3FBE 16'h4740
`define CUBE_LUT_3FBF 16'h4743
`define CUBE_LUT_3FC0 16'h4746
`define CUBE_LUT_3FC1 16'h4749
`define CUBE_LUT_3FC2 16'h474C
`define CUBE_LUT_3FC3 16'h474E
`define CUBE_LUT_3FC4 16'h4751
`define CUBE_LUT_3FC5 16'h4754
`define CUBE_LUT_3FC6 16'h4757
`define CUBE_LUT_3FC7 16'h475A
`define CUBE_LUT_3FC8 16'h475D
`define CUBE_LUT_3FC9 16'h475F
`define CUBE_LUT_3FCA 16'h4762
`define CUBE_LUT_3FCB 16'h4765
`define CUBE_LUT_3FCC 16'h4768
`define CUBE_LUT_3FCD 16'h476B
`define CUBE_LUT_3FCE 16'h476E
`define CUBE_LUT_3FCF 16'h4770
`define CUBE_LUT_3FD0 16'h4773
`define CUBE_LUT_3FD1 16'h4776
`define CUBE_LUT_3FD2 16'h4779
`define CUBE_LUT_3FD3 16'h477C
`define CUBE_LUT_3FD4 16'h477F
`define CUBE_LUT_3FD5 16'h4782
`define CUBE_LUT_3FD6 16'h4785
`define CUBE_LUT_3FD7 16'h4787
`define CUBE_LUT_3FD8 16'h478A
`define CUBE_LUT_3FD9 16'h478D
`define CUBE_LUT_3FDA 16'h4790
`define CUBE_LUT_3FDB 16'h4793
`define CUBE_LUT_3FDC 16'h4796
`define CUBE_LUT_3FDD 16'h4799
`define CUBE_LUT_3FDE 16'h479C
`define CUBE_LUT_3FDF 16'h479F
`define CUBE_LUT_3FE0 16'h47A1
`define CUBE_LUT_3FE1 16'h47A4
`define CUBE_LUT_3FE2 16'h47A7
`define CUBE_LUT_3FE3 16'h47AA
`define CUBE_LUT_3FE4 16'h47AD
`define CUBE_LUT_3FE5 16'h47B0
`define CUBE_LUT_3FE6 16'h47B3
`define CUBE_LUT_3FE7 16'h47B6
`define CUBE_LUT_3FE8 16'h47B9
`define CUBE_LUT_3FE9 16'h47BC
`define CUBE_LUT_3FEA 16'h47BF
`define CUBE_LUT_3FEB 16'h47C2
`define CUBE_LUT_3FEC 16'h47C5
`define CUBE_LUT_3FED 16'h47C8
`define CUBE_LUT_3FEE 16'h47CA
`define CUBE_LUT_3FEF 16'h47CD
`define CUBE_LUT_3FF0 16'h47D0
`define CUBE_LUT_3FF1 16'h47D3
`define CUBE_LUT_3FF2 16'h47D6
`define CUBE_LUT_3FF3 16'h47D9
`define CUBE_LUT_3FF4 16'h47DC
`define CUBE_LUT_3FF5 16'h47DF
`define CUBE_LUT_3FF6 16'h47E2
`define CUBE_LUT_3FF7 16'h47E5
`define CUBE_LUT_3FF8 16'h47E8
`define CUBE_LUT_3FF9 16'h47EB
`define CUBE_LUT_3FFA 16'h47EE
`define CUBE_LUT_3FFB 16'h47F1
`define CUBE_LUT_3FFC 16'h47F4
`define CUBE_LUT_3FFD 16'h47F7
`define CUBE_LUT_3FFE 16'h47FA
`define CUBE_LUT_3FFF 16'h47FD
`define CUBE_LUT_4000 16'h4800
`define CUBE_LUT_4001 16'h4803
`define CUBE_LUT_4002 16'h4806
`define CUBE_LUT_4003 16'h4809
`define CUBE_LUT_4004 16'h480C
`define CUBE_LUT_4005 16'h480F
`define CUBE_LUT_4006 16'h4812
`define CUBE_LUT_4007 16'h4815
`define CUBE_LUT_4008 16'h4818
`define CUBE_LUT_4009 16'h481B
`define CUBE_LUT_400A 16'h481E
`define CUBE_LUT_400B 16'h4821
`define CUBE_LUT_400C 16'h4824
`define CUBE_LUT_400D 16'h4827
`define CUBE_LUT_400E 16'h482B
`define CUBE_LUT_400F 16'h482E
`define CUBE_LUT_4010 16'h4831
`define CUBE_LUT_4011 16'h4834
`define CUBE_LUT_4012 16'h4837
`define CUBE_LUT_4013 16'h483A
`define CUBE_LUT_4014 16'h483D
`define CUBE_LUT_4015 16'h4840
`define CUBE_LUT_4016 16'h4843
`define CUBE_LUT_4017 16'h4847
`define CUBE_LUT_4018 16'h484A
`define CUBE_LUT_4019 16'h484D
`define CUBE_LUT_401A 16'h4850
`define CUBE_LUT_401B 16'h4853
`define CUBE_LUT_401C 16'h4856
`define CUBE_LUT_401D 16'h4859
`define CUBE_LUT_401E 16'h485D
`define CUBE_LUT_401F 16'h4860
`define CUBE_LUT_4020 16'h4863
`define CUBE_LUT_4021 16'h4866
`define CUBE_LUT_4022 16'h4869
`define CUBE_LUT_4023 16'h486D
`define CUBE_LUT_4024 16'h4870
`define CUBE_LUT_4025 16'h4873
`define CUBE_LUT_4026 16'h4876
`define CUBE_LUT_4027 16'h487A
`define CUBE_LUT_4028 16'h487D
`define CUBE_LUT_4029 16'h4880
`define CUBE_LUT_402A 16'h4883
`define CUBE_LUT_402B 16'h4886
`define CUBE_LUT_402C 16'h488A
`define CUBE_LUT_402D 16'h488D
`define CUBE_LUT_402E 16'h4890
`define CUBE_LUT_402F 16'h4894
`define CUBE_LUT_4030 16'h4897
`define CUBE_LUT_4031 16'h489A
`define CUBE_LUT_4032 16'h489D
`define CUBE_LUT_4033 16'h48A1
`define CUBE_LUT_4034 16'h48A4
`define CUBE_LUT_4035 16'h48A7
`define CUBE_LUT_4036 16'h48AB
`define CUBE_LUT_4037 16'h48AE
`define CUBE_LUT_4038 16'h48B1
`define CUBE_LUT_4039 16'h48B5
`define CUBE_LUT_403A 16'h48B8
`define CUBE_LUT_403B 16'h48BB
`define CUBE_LUT_403C 16'h48BF
`define CUBE_LUT_403D 16'h48C2
`define CUBE_LUT_403E 16'h48C5
`define CUBE_LUT_403F 16'h48C9
`define CUBE_LUT_4040 16'h48CC
`define CUBE_LUT_4041 16'h48D0
`define CUBE_LUT_4042 16'h48D3
`define CUBE_LUT_4043 16'h48D6
`define CUBE_LUT_4044 16'h48DA
`define CUBE_LUT_4045 16'h48DD
`define CUBE_LUT_4046 16'h48E1
`define CUBE_LUT_4047 16'h48E4
`define CUBE_LUT_4048 16'h48E8
`define CUBE_LUT_4049 16'h48EB
`define CUBE_LUT_404A 16'h48EE
`define CUBE_LUT_404B 16'h48F2
`define CUBE_LUT_404C 16'h48F5
`define CUBE_LUT_404D 16'h48F9
`define CUBE_LUT_404E 16'h48FC
`define CUBE_LUT_404F 16'h4900
`define CUBE_LUT_4050 16'h4903
`define CUBE_LUT_4051 16'h4907
`define CUBE_LUT_4052 16'h490A
`define CUBE_LUT_4053 16'h490E
`define CUBE_LUT_4054 16'h4911
`define CUBE_LUT_4055 16'h4915
`define CUBE_LUT_4056 16'h4918
`define CUBE_LUT_4057 16'h491C
`define CUBE_LUT_4058 16'h491F
`define CUBE_LUT_4059 16'h4923
`define CUBE_LUT_405A 16'h4926
`define CUBE_LUT_405B 16'h492A
`define CUBE_LUT_405C 16'h492E
`define CUBE_LUT_405D 16'h4931
`define CUBE_LUT_405E 16'h4935
`define CUBE_LUT_405F 16'h4938
`define CUBE_LUT_4060 16'h493C
`define CUBE_LUT_4061 16'h493F
`define CUBE_LUT_4062 16'h4943
`define CUBE_LUT_4063 16'h4947
`define CUBE_LUT_4064 16'h494A
`define CUBE_LUT_4065 16'h494E
`define CUBE_LUT_4066 16'h4951
`define CUBE_LUT_4067 16'h4955
`define CUBE_LUT_4068 16'h4959
`define CUBE_LUT_4069 16'h495C
`define CUBE_LUT_406A 16'h4960
`define CUBE_LUT_406B 16'h4964
`define CUBE_LUT_406C 16'h4967
`define CUBE_LUT_406D 16'h496B
`define CUBE_LUT_406E 16'h496F
`define CUBE_LUT_406F 16'h4972
`define CUBE_LUT_4070 16'h4976
`define CUBE_LUT_4071 16'h497A
`define CUBE_LUT_4072 16'h497D
`define CUBE_LUT_4073 16'h4981
`define CUBE_LUT_4074 16'h4985
`define CUBE_LUT_4075 16'h4989
`define CUBE_LUT_4076 16'h498C
`define CUBE_LUT_4077 16'h4990
`define CUBE_LUT_4078 16'h4994
`define CUBE_LUT_4079 16'h4998
`define CUBE_LUT_407A 16'h499B
`define CUBE_LUT_407B 16'h499F
`define CUBE_LUT_407C 16'h49A3
`define CUBE_LUT_407D 16'h49A7
`define CUBE_LUT_407E 16'h49AA
`define CUBE_LUT_407F 16'h49AE
`define CUBE_LUT_4080 16'h49B2
`define CUBE_LUT_4081 16'h49B6
`define CUBE_LUT_4082 16'h49BA
`define CUBE_LUT_4083 16'h49BD
`define CUBE_LUT_4084 16'h49C1
`define CUBE_LUT_4085 16'h49C5
`define CUBE_LUT_4086 16'h49C9
`define CUBE_LUT_4087 16'h49CD
`define CUBE_LUT_4088 16'h49D1
`define CUBE_LUT_4089 16'h49D4
`define CUBE_LUT_408A 16'h49D8
`define CUBE_LUT_408B 16'h49DC
`define CUBE_LUT_408C 16'h49E0
`define CUBE_LUT_408D 16'h49E4
`define CUBE_LUT_408E 16'h49E8
`define CUBE_LUT_408F 16'h49EC
`define CUBE_LUT_4090 16'h49F0
`define CUBE_LUT_4091 16'h49F4
`define CUBE_LUT_4092 16'h49F7
`define CUBE_LUT_4093 16'h49FB
`define CUBE_LUT_4094 16'h49FF
`define CUBE_LUT_4095 16'h4A03
`define CUBE_LUT_4096 16'h4A07
`define CUBE_LUT_4097 16'h4A0B
`define CUBE_LUT_4098 16'h4A0F
`define CUBE_LUT_4099 16'h4A13
`define CUBE_LUT_409A 16'h4A17
`define CUBE_LUT_409B 16'h4A1B
`define CUBE_LUT_409C 16'h4A1F
`define CUBE_LUT_409D 16'h4A23
`define CUBE_LUT_409E 16'h4A27
`define CUBE_LUT_409F 16'h4A2B
`define CUBE_LUT_40A0 16'h4A2F
`define CUBE_LUT_40A1 16'h4A33
`define CUBE_LUT_40A2 16'h4A37
`define CUBE_LUT_40A3 16'h4A3B
`define CUBE_LUT_40A4 16'h4A3F
`define CUBE_LUT_40A5 16'h4A43
`define CUBE_LUT_40A6 16'h4A47
`define CUBE_LUT_40A7 16'h4A4B
`define CUBE_LUT_40A8 16'h4A4F
`define CUBE_LUT_40A9 16'h4A53
`define CUBE_LUT_40AA 16'h4A57
`define CUBE_LUT_40AB 16'h4A5B
`define CUBE_LUT_40AC 16'h4A60
`define CUBE_LUT_40AD 16'h4A64
`define CUBE_LUT_40AE 16'h4A68
`define CUBE_LUT_40AF 16'h4A6C
`define CUBE_LUT_40B0 16'h4A70
`define CUBE_LUT_40B1 16'h4A74
`define CUBE_LUT_40B2 16'h4A78
`define CUBE_LUT_40B3 16'h4A7C
`define CUBE_LUT_40B4 16'h4A80
`define CUBE_LUT_40B5 16'h4A85
`define CUBE_LUT_40B6 16'h4A89
`define CUBE_LUT_40B7 16'h4A8D
`define CUBE_LUT_40B8 16'h4A91
`define CUBE_LUT_40B9 16'h4A95
`define CUBE_LUT_40BA 16'h4A99
`define CUBE_LUT_40BB 16'h4A9E
`define CUBE_LUT_40BC 16'h4AA2
`define CUBE_LUT_40BD 16'h4AA6
`define CUBE_LUT_40BE 16'h4AAA
`define CUBE_LUT_40BF 16'h4AAF
`define CUBE_LUT_40C0 16'h4AB3
`define CUBE_LUT_40C1 16'h4AB7
`define CUBE_LUT_40C2 16'h4ABB
`define CUBE_LUT_40C3 16'h4ABF
`define CUBE_LUT_40C4 16'h4AC4
`define CUBE_LUT_40C5 16'h4AC8
`define CUBE_LUT_40C6 16'h4ACC
`define CUBE_LUT_40C7 16'h4AD1
`define CUBE_LUT_40C8 16'h4AD5
`define CUBE_LUT_40C9 16'h4AD9
`define CUBE_LUT_40CA 16'h4ADD
`define CUBE_LUT_40CB 16'h4AE2
`define CUBE_LUT_40CC 16'h4AE6
`define CUBE_LUT_40CD 16'h4AEA
`define CUBE_LUT_40CE 16'h4AEF
`define CUBE_LUT_40CF 16'h4AF3
`define CUBE_LUT_40D0 16'h4AF7
`define CUBE_LUT_40D1 16'h4AFC
`define CUBE_LUT_40D2 16'h4B00
`define CUBE_LUT_40D3 16'h4B04
`define CUBE_LUT_40D4 16'h4B09
`define CUBE_LUT_40D5 16'h4B0D
`define CUBE_LUT_40D6 16'h4B12
`define CUBE_LUT_40D7 16'h4B16
`define CUBE_LUT_40D8 16'h4B1A
`define CUBE_LUT_40D9 16'h4B1F
`define CUBE_LUT_40DA 16'h4B23
`define CUBE_LUT_40DB 16'h4B28
`define CUBE_LUT_40DC 16'h4B2C
`define CUBE_LUT_40DD 16'h4B30
`define CUBE_LUT_40DE 16'h4B35
`define CUBE_LUT_40DF 16'h4B39
`define CUBE_LUT_40E0 16'h4B3E
`define CUBE_LUT_40E1 16'h4B42
`define CUBE_LUT_40E2 16'h4B47
`define CUBE_LUT_40E3 16'h4B4B
`define CUBE_LUT_40E4 16'h4B50
`define CUBE_LUT_40E5 16'h4B54
`define CUBE_LUT_40E6 16'h4B59
`define CUBE_LUT_40E7 16'h4B5D
`define CUBE_LUT_40E8 16'h4B62
`define CUBE_LUT_40E9 16'h4B66
`define CUBE_LUT_40EA 16'h4B6B
`define CUBE_LUT_40EB 16'h4B6F
`define CUBE_LUT_40EC 16'h4B74
`define CUBE_LUT_40ED 16'h4B78
`define CUBE_LUT_40EE 16'h4B7D
`define CUBE_LUT_40EF 16'h4B81
`define CUBE_LUT_40F0 16'h4B86
`define CUBE_LUT_40F1 16'h4B8B
`define CUBE_LUT_40F2 16'h4B8F
`define CUBE_LUT_40F3 16'h4B94
`define CUBE_LUT_40F4 16'h4B98
`define CUBE_LUT_40F5 16'h4B9D
`define CUBE_LUT_40F6 16'h4BA1
`define CUBE_LUT_40F7 16'h4BA6
`define CUBE_LUT_40F8 16'h4BAB
`define CUBE_LUT_40F9 16'h4BAF
`define CUBE_LUT_40FA 16'h4BB4
`define CUBE_LUT_40FB 16'h4BB9
`define CUBE_LUT_40FC 16'h4BBD
`define CUBE_LUT_40FD 16'h4BC2
`define CUBE_LUT_40FE 16'h4BC7
`define CUBE_LUT_40FF 16'h4BCB
`define CUBE_LUT_4100 16'h4BD0
`define CUBE_LUT_4101 16'h4BD5
`define CUBE_LUT_4102 16'h4BD9
`define CUBE_LUT_4103 16'h4BDE
`define CUBE_LUT_4104 16'h4BE3
`define CUBE_LUT_4105 16'h4BE8
`define CUBE_LUT_4106 16'h4BEC
`define CUBE_LUT_4107 16'h4BF1
`define CUBE_LUT_4108 16'h4BF6
`define CUBE_LUT_4109 16'h4BFA
`define CUBE_LUT_410A 16'h4BFF
`define CUBE_LUT_410B 16'h4C02
`define CUBE_LUT_410C 16'h4C04
`define CUBE_LUT_410D 16'h4C07
`define CUBE_LUT_410E 16'h4C09
`define CUBE_LUT_410F 16'h4C0C
`define CUBE_LUT_4110 16'h4C0E
`define CUBE_LUT_4111 16'h4C10
`define CUBE_LUT_4112 16'h4C13
`define CUBE_LUT_4113 16'h4C15
`define CUBE_LUT_4114 16'h4C18
`define CUBE_LUT_4115 16'h4C1A
`define CUBE_LUT_4116 16'h4C1C
`define CUBE_LUT_4117 16'h4C1F
`define CUBE_LUT_4118 16'h4C21
`define CUBE_LUT_4119 16'h4C24
`define CUBE_LUT_411A 16'h4C26
`define CUBE_LUT_411B 16'h4C29
`define CUBE_LUT_411C 16'h4C2B
`define CUBE_LUT_411D 16'h4C2E
`define CUBE_LUT_411E 16'h4C30
`define CUBE_LUT_411F 16'h4C32
`define CUBE_LUT_4120 16'h4C35
`define CUBE_LUT_4121 16'h4C37
`define CUBE_LUT_4122 16'h4C3A
`define CUBE_LUT_4123 16'h4C3C
`define CUBE_LUT_4124 16'h4C3F
`define CUBE_LUT_4125 16'h4C41
`define CUBE_LUT_4126 16'h4C44
`define CUBE_LUT_4127 16'h4C46
`define CUBE_LUT_4128 16'h4C49
`define CUBE_LUT_4129 16'h4C4B
`define CUBE_LUT_412A 16'h4C4E
`define CUBE_LUT_412B 16'h4C50
`define CUBE_LUT_412C 16'h4C53
`define CUBE_LUT_412D 16'h4C55
`define CUBE_LUT_412E 16'h4C58
`define CUBE_LUT_412F 16'h4C5A
`define CUBE_LUT_4130 16'h4C5D
`define CUBE_LUT_4131 16'h4C5F
`define CUBE_LUT_4132 16'h4C62
`define CUBE_LUT_4133 16'h4C64
`define CUBE_LUT_4134 16'h4C67
`define CUBE_LUT_4135 16'h4C69
`define CUBE_LUT_4136 16'h4C6C
`define CUBE_LUT_4137 16'h4C6F
`define CUBE_LUT_4138 16'h4C71
`define CUBE_LUT_4139 16'h4C74
`define CUBE_LUT_413A 16'h4C76
`define CUBE_LUT_413B 16'h4C79
`define CUBE_LUT_413C 16'h4C7B
`define CUBE_LUT_413D 16'h4C7E
`define CUBE_LUT_413E 16'h4C80
`define CUBE_LUT_413F 16'h4C83
`define CUBE_LUT_4140 16'h4C86
`define CUBE_LUT_4141 16'h4C88
`define CUBE_LUT_4142 16'h4C8B
`define CUBE_LUT_4143 16'h4C8D
`define CUBE_LUT_4144 16'h4C90
`define CUBE_LUT_4145 16'h4C93
`define CUBE_LUT_4146 16'h4C95
`define CUBE_LUT_4147 16'h4C98
`define CUBE_LUT_4148 16'h4C9A
`define CUBE_LUT_4149 16'h4C9D
`define CUBE_LUT_414A 16'h4CA0
`define CUBE_LUT_414B 16'h4CA2
`define CUBE_LUT_414C 16'h4CA5
`define CUBE_LUT_414D 16'h4CA8
`define CUBE_LUT_414E 16'h4CAA
`define CUBE_LUT_414F 16'h4CAD
`define CUBE_LUT_4150 16'h4CAF
`define CUBE_LUT_4151 16'h4CB2
`define CUBE_LUT_4152 16'h4CB5
`define CUBE_LUT_4153 16'h4CB7
`define CUBE_LUT_4154 16'h4CBA
`define CUBE_LUT_4155 16'h4CBD
`define CUBE_LUT_4156 16'h4CBF
`define CUBE_LUT_4157 16'h4CC2
`define CUBE_LUT_4158 16'h4CC5
`define CUBE_LUT_4159 16'h4CC7
`define CUBE_LUT_415A 16'h4CCA
`define CUBE_LUT_415B 16'h4CCD
`define CUBE_LUT_415C 16'h4CCF
`define CUBE_LUT_415D 16'h4CD2
`define CUBE_LUT_415E 16'h4CD5
`define CUBE_LUT_415F 16'h4CD8
`define CUBE_LUT_4160 16'h4CDA
`define CUBE_LUT_4161 16'h4CDD
`define CUBE_LUT_4162 16'h4CE0
`define CUBE_LUT_4163 16'h4CE2
`define CUBE_LUT_4164 16'h4CE5
`define CUBE_LUT_4165 16'h4CE8
`define CUBE_LUT_4166 16'h4CEB
`define CUBE_LUT_4167 16'h4CED
`define CUBE_LUT_4168 16'h4CF0
`define CUBE_LUT_4169 16'h4CF3
`define CUBE_LUT_416A 16'h4CF6
`define CUBE_LUT_416B 16'h4CF8
`define CUBE_LUT_416C 16'h4CFB
`define CUBE_LUT_416D 16'h4CFE
`define CUBE_LUT_416E 16'h4D01
`define CUBE_LUT_416F 16'h4D03
`define CUBE_LUT_4170 16'h4D06
`define CUBE_LUT_4171 16'h4D09
`define CUBE_LUT_4172 16'h4D0C
`define CUBE_LUT_4173 16'h4D0E
`define CUBE_LUT_4174 16'h4D11
`define CUBE_LUT_4175 16'h4D14
`define CUBE_LUT_4176 16'h4D17
`define CUBE_LUT_4177 16'h4D1A
`define CUBE_LUT_4178 16'h4D1C
`define CUBE_LUT_4179 16'h4D1F
`define CUBE_LUT_417A 16'h4D22
`define CUBE_LUT_417B 16'h4D25
`define CUBE_LUT_417C 16'h4D28
`define CUBE_LUT_417D 16'h4D2B
`define CUBE_LUT_417E 16'h4D2D
`define CUBE_LUT_417F 16'h4D30
`define CUBE_LUT_4180 16'h4D33
`define CUBE_LUT_4181 16'h4D36
`define CUBE_LUT_4182 16'h4D39
`define CUBE_LUT_4183 16'h4D3C
`define CUBE_LUT_4184 16'h4D3E
`define CUBE_LUT_4185 16'h4D41
`define CUBE_LUT_4186 16'h4D44
`define CUBE_LUT_4187 16'h4D47
`define CUBE_LUT_4188 16'h4D4A
`define CUBE_LUT_4189 16'h4D4D
`define CUBE_LUT_418A 16'h4D50
`define CUBE_LUT_418B 16'h4D52
`define CUBE_LUT_418C 16'h4D55
`define CUBE_LUT_418D 16'h4D58
`define CUBE_LUT_418E 16'h4D5B
`define CUBE_LUT_418F 16'h4D5E
`define CUBE_LUT_4190 16'h4D61
`define CUBE_LUT_4191 16'h4D64
`define CUBE_LUT_4192 16'h4D67
`define CUBE_LUT_4193 16'h4D6A
`define CUBE_LUT_4194 16'h4D6D
`define CUBE_LUT_4195 16'h4D6F
`define CUBE_LUT_4196 16'h4D72
`define CUBE_LUT_4197 16'h4D75
`define CUBE_LUT_4198 16'h4D78
`define CUBE_LUT_4199 16'h4D7B
`define CUBE_LUT_419A 16'h4D7E
`define CUBE_LUT_419B 16'h4D81
`define CUBE_LUT_419C 16'h4D84
`define CUBE_LUT_419D 16'h4D87
`define CUBE_LUT_419E 16'h4D8A
`define CUBE_LUT_419F 16'h4D8D
`define CUBE_LUT_41A0 16'h4D90
`define CUBE_LUT_41A1 16'h4D93
`define CUBE_LUT_41A2 16'h4D96
`define CUBE_LUT_41A3 16'h4D99
`define CUBE_LUT_41A4 16'h4D9C
`define CUBE_LUT_41A5 16'h4D9F
`define CUBE_LUT_41A6 16'h4DA2
`define CUBE_LUT_41A7 16'h4DA5
`define CUBE_LUT_41A8 16'h4DA8
`define CUBE_LUT_41A9 16'h4DAB
`define CUBE_LUT_41AA 16'h4DAE
`define CUBE_LUT_41AB 16'h4DB1
`define CUBE_LUT_41AC 16'h4DB4
`define CUBE_LUT_41AD 16'h4DB7
`define CUBE_LUT_41AE 16'h4DBA
`define CUBE_LUT_41AF 16'h4DBD
`define CUBE_LUT_41B0 16'h4DC0
`define CUBE_LUT_41B1 16'h4DC3
`define CUBE_LUT_41B2 16'h4DC6
`define CUBE_LUT_41B3 16'h4DC9
`define CUBE_LUT_41B4 16'h4DCC
`define CUBE_LUT_41B5 16'h4DCF
`define CUBE_LUT_41B6 16'h4DD2
`define CUBE_LUT_41B7 16'h4DD5
`define CUBE_LUT_41B8 16'h4DD8
`define CUBE_LUT_41B9 16'h4DDB
`define CUBE_LUT_41BA 16'h4DDE
`define CUBE_LUT_41BB 16'h4DE1
`define CUBE_LUT_41BC 16'h4DE5
`define CUBE_LUT_41BD 16'h4DE8
`define CUBE_LUT_41BE 16'h4DEB
`define CUBE_LUT_41BF 16'h4DEE
`define CUBE_LUT_41C0 16'h4DF1
`define CUBE_LUT_41C1 16'h4DF4
`define CUBE_LUT_41C2 16'h4DF7
`define CUBE_LUT_41C3 16'h4DFA
`define CUBE_LUT_41C4 16'h4DFD
`define CUBE_LUT_41C5 16'h4E00
`define CUBE_LUT_41C6 16'h4E04
`define CUBE_LUT_41C7 16'h4E07
`define CUBE_LUT_41C8 16'h4E0A
`define CUBE_LUT_41C9 16'h4E0D
`define CUBE_LUT_41CA 16'h4E10
`define CUBE_LUT_41CB 16'h4E13
`define CUBE_LUT_41CC 16'h4E16
`define CUBE_LUT_41CD 16'h4E1A
`define CUBE_LUT_41CE 16'h4E1D
`define CUBE_LUT_41CF 16'h4E20
`define CUBE_LUT_41D0 16'h4E23
`define CUBE_LUT_41D1 16'h4E26
`define CUBE_LUT_41D2 16'h4E29
`define CUBE_LUT_41D3 16'h4E2D
`define CUBE_LUT_41D4 16'h4E30
`define CUBE_LUT_41D5 16'h4E33
`define CUBE_LUT_41D6 16'h4E36
`define CUBE_LUT_41D7 16'h4E39
`define CUBE_LUT_41D8 16'h4E3C
`define CUBE_LUT_41D9 16'h4E40
`define CUBE_LUT_41DA 16'h4E43
`define CUBE_LUT_41DB 16'h4E46
`define CUBE_LUT_41DC 16'h4E49
`define CUBE_LUT_41DD 16'h4E4D
`define CUBE_LUT_41DE 16'h4E50
`define CUBE_LUT_41DF 16'h4E53
`define CUBE_LUT_41E0 16'h4E56
`define CUBE_LUT_41E1 16'h4E59
`define CUBE_LUT_41E2 16'h4E5D
`define CUBE_LUT_41E3 16'h4E60
`define CUBE_LUT_41E4 16'h4E63
`define CUBE_LUT_41E5 16'h4E66
`define CUBE_LUT_41E6 16'h4E6A
`define CUBE_LUT_41E7 16'h4E6D
`define CUBE_LUT_41E8 16'h4E70
`define CUBE_LUT_41E9 16'h4E74
`define CUBE_LUT_41EA 16'h4E77
`define CUBE_LUT_41EB 16'h4E7A
`define CUBE_LUT_41EC 16'h4E7D
`define CUBE_LUT_41ED 16'h4E81
`define CUBE_LUT_41EE 16'h4E84
`define CUBE_LUT_41EF 16'h4E87
`define CUBE_LUT_41F0 16'h4E8B
`define CUBE_LUT_41F1 16'h4E8E
`define CUBE_LUT_41F2 16'h4E91
`define CUBE_LUT_41F3 16'h4E94
`define CUBE_LUT_41F4 16'h4E98
`define CUBE_LUT_41F5 16'h4E9B
`define CUBE_LUT_41F6 16'h4E9E
`define CUBE_LUT_41F7 16'h4EA2
`define CUBE_LUT_41F8 16'h4EA5
`define CUBE_LUT_41F9 16'h4EA8
`define CUBE_LUT_41FA 16'h4EAC
`define CUBE_LUT_41FB 16'h4EAF
`define CUBE_LUT_41FC 16'h4EB3
`define CUBE_LUT_41FD 16'h4EB6
`define CUBE_LUT_41FE 16'h4EB9
`define CUBE_LUT_41FF 16'h4EBD
`define CUBE_LUT_4200 16'h4EC0
