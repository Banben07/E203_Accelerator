`define TANH_LUT_NEGATIVE_SIZE 2140
`define TANH_LUT_NEGATIVE_BITS 12
`define TANH_LUT_NEGATIVE_8000 16'h8000
`define TANH_LUT_NEGATIVE_8008 16'h8008
`define TANH_LUT_NEGATIVE_8010 16'h8010
`define TANH_LUT_NEGATIVE_8018 16'h8018
`define TANH_LUT_NEGATIVE_8020 16'h8020
`define TANH_LUT_NEGATIVE_8028 16'h8028
`define TANH_LUT_NEGATIVE_8030 16'h8030
`define TANH_LUT_NEGATIVE_8038 16'h8038
`define TANH_LUT_NEGATIVE_8040 16'h8040
`define TANH_LUT_NEGATIVE_8048 16'h8048
`define TANH_LUT_NEGATIVE_8050 16'h8050
`define TANH_LUT_NEGATIVE_8058 16'h8058
`define TANH_LUT_NEGATIVE_8060 16'h8060
`define TANH_LUT_NEGATIVE_8068 16'h8068
`define TANH_LUT_NEGATIVE_8070 16'h8070
`define TANH_LUT_NEGATIVE_8078 16'h8078
`define TANH_LUT_NEGATIVE_8080 16'h8080
`define TANH_LUT_NEGATIVE_8088 16'h8088
`define TANH_LUT_NEGATIVE_8090 16'h8090
`define TANH_LUT_NEGATIVE_8098 16'h8098
`define TANH_LUT_NEGATIVE_80A0 16'h80A0
`define TANH_LUT_NEGATIVE_80A8 16'h80A8
`define TANH_LUT_NEGATIVE_80B0 16'h80B0
`define TANH_LUT_NEGATIVE_80B8 16'h80B8
`define TANH_LUT_NEGATIVE_80C0 16'h80C0
`define TANH_LUT_NEGATIVE_80C8 16'h80C8
`define TANH_LUT_NEGATIVE_80D0 16'h80D0
`define TANH_LUT_NEGATIVE_80D8 16'h80D8
`define TANH_LUT_NEGATIVE_80E0 16'h80E0
`define TANH_LUT_NEGATIVE_80E8 16'h80E8
`define TANH_LUT_NEGATIVE_80F0 16'h80F0
`define TANH_LUT_NEGATIVE_80F8 16'h80F8
`define TANH_LUT_NEGATIVE_8100 16'h8100
`define TANH_LUT_NEGATIVE_8108 16'h8108
`define TANH_LUT_NEGATIVE_8110 16'h8110
`define TANH_LUT_NEGATIVE_8118 16'h8118
`define TANH_LUT_NEGATIVE_8120 16'h8120
`define TANH_LUT_NEGATIVE_8128 16'h8128
`define TANH_LUT_NEGATIVE_8130 16'h8130
`define TANH_LUT_NEGATIVE_8138 16'h8138
`define TANH_LUT_NEGATIVE_8140 16'h8140
`define TANH_LUT_NEGATIVE_8148 16'h8148
`define TANH_LUT_NEGATIVE_8150 16'h8150
`define TANH_LUT_NEGATIVE_8158 16'h8158
`define TANH_LUT_NEGATIVE_8160 16'h8160
`define TANH_LUT_NEGATIVE_8168 16'h8168
`define TANH_LUT_NEGATIVE_8170 16'h8170
`define TANH_LUT_NEGATIVE_8178 16'h8178
`define TANH_LUT_NEGATIVE_8180 16'h8180
`define TANH_LUT_NEGATIVE_8188 16'h8188
`define TANH_LUT_NEGATIVE_8190 16'h8190
`define TANH_LUT_NEGATIVE_8198 16'h8198
`define TANH_LUT_NEGATIVE_81A0 16'h81A0
`define TANH_LUT_NEGATIVE_81A8 16'h81A8
`define TANH_LUT_NEGATIVE_81B0 16'h81B0
`define TANH_LUT_NEGATIVE_81B8 16'h81B8
`define TANH_LUT_NEGATIVE_81C0 16'h81C0
`define TANH_LUT_NEGATIVE_81C8 16'h81C8
`define TANH_LUT_NEGATIVE_81D0 16'h81D0
`define TANH_LUT_NEGATIVE_81D8 16'h81D8
`define TANH_LUT_NEGATIVE_81E0 16'h81E0
`define TANH_LUT_NEGATIVE_81E8 16'h81E8
`define TANH_LUT_NEGATIVE_81F0 16'h81F0
`define TANH_LUT_NEGATIVE_81F8 16'h81F8
`define TANH_LUT_NEGATIVE_8200 16'h8200
`define TANH_LUT_NEGATIVE_8208 16'h8208
`define TANH_LUT_NEGATIVE_8210 16'h8210
`define TANH_LUT_NEGATIVE_8218 16'h8218
`define TANH_LUT_NEGATIVE_8220 16'h8220
`define TANH_LUT_NEGATIVE_8228 16'h8228
`define TANH_LUT_NEGATIVE_8230 16'h8230
`define TANH_LUT_NEGATIVE_8238 16'h8238
`define TANH_LUT_NEGATIVE_8240 16'h8240
`define TANH_LUT_NEGATIVE_8248 16'h8248
`define TANH_LUT_NEGATIVE_8250 16'h8250
`define TANH_LUT_NEGATIVE_8258 16'h8258
`define TANH_LUT_NEGATIVE_8260 16'h8260
`define TANH_LUT_NEGATIVE_8268 16'h8268
`define TANH_LUT_NEGATIVE_8270 16'h8270
`define TANH_LUT_NEGATIVE_8278 16'h8278
`define TANH_LUT_NEGATIVE_8280 16'h8280
`define TANH_LUT_NEGATIVE_8288 16'h8288
`define TANH_LUT_NEGATIVE_8290 16'h8290
`define TANH_LUT_NEGATIVE_8298 16'h8298
`define TANH_LUT_NEGATIVE_82A0 16'h82A0
`define TANH_LUT_NEGATIVE_82A8 16'h82A8
`define TANH_LUT_NEGATIVE_82B0 16'h82B0
`define TANH_LUT_NEGATIVE_82B8 16'h82B8
`define TANH_LUT_NEGATIVE_82C0 16'h82C0
`define TANH_LUT_NEGATIVE_82C8 16'h82C8
`define TANH_LUT_NEGATIVE_82D0 16'h82D0
`define TANH_LUT_NEGATIVE_82D8 16'h82D8
`define TANH_LUT_NEGATIVE_82E0 16'h82E0
`define TANH_LUT_NEGATIVE_82E8 16'h82E8
`define TANH_LUT_NEGATIVE_82F0 16'h82F0
`define TANH_LUT_NEGATIVE_82F8 16'h82F8
`define TANH_LUT_NEGATIVE_8300 16'h8300
`define TANH_LUT_NEGATIVE_8308 16'h8308
`define TANH_LUT_NEGATIVE_8310 16'h8310
`define TANH_LUT_NEGATIVE_8318 16'h8318
`define TANH_LUT_NEGATIVE_8320 16'h8320
`define TANH_LUT_NEGATIVE_8328 16'h8328
`define TANH_LUT_NEGATIVE_8330 16'h8330
`define TANH_LUT_NEGATIVE_8338 16'h8338
`define TANH_LUT_NEGATIVE_8340 16'h8340
`define TANH_LUT_NEGATIVE_8348 16'h8348
`define TANH_LUT_NEGATIVE_8350 16'h8350
`define TANH_LUT_NEGATIVE_8358 16'h8358
`define TANH_LUT_NEGATIVE_8360 16'h8360
`define TANH_LUT_NEGATIVE_8368 16'h8368
`define TANH_LUT_NEGATIVE_8370 16'h8370
`define TANH_LUT_NEGATIVE_8378 16'h8378
`define TANH_LUT_NEGATIVE_8380 16'h8380
`define TANH_LUT_NEGATIVE_8388 16'h8388
`define TANH_LUT_NEGATIVE_8390 16'h8390
`define TANH_LUT_NEGATIVE_8398 16'h8398
`define TANH_LUT_NEGATIVE_83A0 16'h83A0
`define TANH_LUT_NEGATIVE_83A8 16'h83A8
`define TANH_LUT_NEGATIVE_83B0 16'h83B0
`define TANH_LUT_NEGATIVE_83B8 16'h83B8
`define TANH_LUT_NEGATIVE_83C0 16'h83C0
`define TANH_LUT_NEGATIVE_83C8 16'h83C8
`define TANH_LUT_NEGATIVE_83D0 16'h83D0
`define TANH_LUT_NEGATIVE_83D8 16'h83D8
`define TANH_LUT_NEGATIVE_83E0 16'h83E0
`define TANH_LUT_NEGATIVE_83E8 16'h83E8
`define TANH_LUT_NEGATIVE_83F0 16'h83F0
`define TANH_LUT_NEGATIVE_83F8 16'h83F8
`define TANH_LUT_NEGATIVE_8400 16'h8400
`define TANH_LUT_NEGATIVE_8408 16'h8408
`define TANH_LUT_NEGATIVE_8410 16'h8410
`define TANH_LUT_NEGATIVE_8418 16'h8418
`define TANH_LUT_NEGATIVE_8420 16'h8420
`define TANH_LUT_NEGATIVE_8428 16'h8428
`define TANH_LUT_NEGATIVE_8430 16'h8430
`define TANH_LUT_NEGATIVE_8438 16'h8438
`define TANH_LUT_NEGATIVE_8440 16'h8440
`define TANH_LUT_NEGATIVE_8448 16'h8448
`define TANH_LUT_NEGATIVE_8450 16'h8450
`define TANH_LUT_NEGATIVE_8458 16'h8458
`define TANH_LUT_NEGATIVE_8460 16'h8460
`define TANH_LUT_NEGATIVE_8468 16'h8468
`define TANH_LUT_NEGATIVE_8470 16'h8470
`define TANH_LUT_NEGATIVE_8478 16'h8478
`define TANH_LUT_NEGATIVE_8480 16'h8480
`define TANH_LUT_NEGATIVE_8488 16'h8488
`define TANH_LUT_NEGATIVE_8490 16'h8490
`define TANH_LUT_NEGATIVE_8498 16'h8498
`define TANH_LUT_NEGATIVE_84A0 16'h84A0
`define TANH_LUT_NEGATIVE_84A8 16'h84A8
`define TANH_LUT_NEGATIVE_84B0 16'h84B0
`define TANH_LUT_NEGATIVE_84B8 16'h84B8
`define TANH_LUT_NEGATIVE_84C0 16'h84C0
`define TANH_LUT_NEGATIVE_84C8 16'h84C8
`define TANH_LUT_NEGATIVE_84D0 16'h84D0
`define TANH_LUT_NEGATIVE_84D8 16'h84D8
`define TANH_LUT_NEGATIVE_84E0 16'h84E0
`define TANH_LUT_NEGATIVE_84E8 16'h84E8
`define TANH_LUT_NEGATIVE_84F0 16'h84F0
`define TANH_LUT_NEGATIVE_84F8 16'h84F8
`define TANH_LUT_NEGATIVE_8500 16'h8500
`define TANH_LUT_NEGATIVE_8508 16'h8508
`define TANH_LUT_NEGATIVE_8510 16'h8510
`define TANH_LUT_NEGATIVE_8518 16'h8518
`define TANH_LUT_NEGATIVE_8520 16'h8520
`define TANH_LUT_NEGATIVE_8528 16'h8528
`define TANH_LUT_NEGATIVE_8530 16'h8530
`define TANH_LUT_NEGATIVE_8538 16'h8538
`define TANH_LUT_NEGATIVE_8540 16'h8540
`define TANH_LUT_NEGATIVE_8548 16'h8548
`define TANH_LUT_NEGATIVE_8550 16'h8550
`define TANH_LUT_NEGATIVE_8558 16'h8558
`define TANH_LUT_NEGATIVE_8560 16'h8560
`define TANH_LUT_NEGATIVE_8568 16'h8568
`define TANH_LUT_NEGATIVE_8570 16'h8570
`define TANH_LUT_NEGATIVE_8578 16'h8578
`define TANH_LUT_NEGATIVE_8580 16'h8580
`define TANH_LUT_NEGATIVE_8588 16'h8588
`define TANH_LUT_NEGATIVE_8590 16'h8590
`define TANH_LUT_NEGATIVE_8598 16'h8598
`define TANH_LUT_NEGATIVE_85A0 16'h85A0
`define TANH_LUT_NEGATIVE_85A8 16'h85A8
`define TANH_LUT_NEGATIVE_85B0 16'h85B0
`define TANH_LUT_NEGATIVE_85B8 16'h85B8
`define TANH_LUT_NEGATIVE_85C0 16'h85C0
`define TANH_LUT_NEGATIVE_85C8 16'h85C8
`define TANH_LUT_NEGATIVE_85D0 16'h85D0
`define TANH_LUT_NEGATIVE_85D8 16'h85D8
`define TANH_LUT_NEGATIVE_85E0 16'h85E0
`define TANH_LUT_NEGATIVE_85E8 16'h85E8
`define TANH_LUT_NEGATIVE_85F0 16'h85F0
`define TANH_LUT_NEGATIVE_85F8 16'h85F8
`define TANH_LUT_NEGATIVE_8600 16'h8600
`define TANH_LUT_NEGATIVE_8608 16'h8608
`define TANH_LUT_NEGATIVE_8610 16'h8610
`define TANH_LUT_NEGATIVE_8618 16'h8618
`define TANH_LUT_NEGATIVE_8620 16'h8620
`define TANH_LUT_NEGATIVE_8628 16'h8628
`define TANH_LUT_NEGATIVE_8630 16'h8630
`define TANH_LUT_NEGATIVE_8638 16'h8638
`define TANH_LUT_NEGATIVE_8640 16'h8640
`define TANH_LUT_NEGATIVE_8648 16'h8648
`define TANH_LUT_NEGATIVE_8650 16'h8650
`define TANH_LUT_NEGATIVE_8658 16'h8658
`define TANH_LUT_NEGATIVE_8660 16'h8660
`define TANH_LUT_NEGATIVE_8668 16'h8668
`define TANH_LUT_NEGATIVE_8670 16'h8670
`define TANH_LUT_NEGATIVE_8678 16'h8678
`define TANH_LUT_NEGATIVE_8680 16'h8680
`define TANH_LUT_NEGATIVE_8688 16'h8688
`define TANH_LUT_NEGATIVE_8690 16'h8690
`define TANH_LUT_NEGATIVE_8698 16'h8698
`define TANH_LUT_NEGATIVE_86A0 16'h86A0
`define TANH_LUT_NEGATIVE_86A8 16'h86A8
`define TANH_LUT_NEGATIVE_86B0 16'h86B0
`define TANH_LUT_NEGATIVE_86B8 16'h86B8
`define TANH_LUT_NEGATIVE_86C0 16'h86C0
`define TANH_LUT_NEGATIVE_86C8 16'h86C8
`define TANH_LUT_NEGATIVE_86D0 16'h86D0
`define TANH_LUT_NEGATIVE_86D8 16'h86D8
`define TANH_LUT_NEGATIVE_86E0 16'h86E0
`define TANH_LUT_NEGATIVE_86E8 16'h86E8
`define TANH_LUT_NEGATIVE_86F0 16'h86F0
`define TANH_LUT_NEGATIVE_86F8 16'h86F8
`define TANH_LUT_NEGATIVE_8700 16'h8700
`define TANH_LUT_NEGATIVE_8708 16'h8708
`define TANH_LUT_NEGATIVE_8710 16'h8710
`define TANH_LUT_NEGATIVE_8718 16'h8718
`define TANH_LUT_NEGATIVE_8720 16'h8720
`define TANH_LUT_NEGATIVE_8728 16'h8728
`define TANH_LUT_NEGATIVE_8730 16'h8730
`define TANH_LUT_NEGATIVE_8738 16'h8738
`define TANH_LUT_NEGATIVE_8740 16'h8740
`define TANH_LUT_NEGATIVE_8748 16'h8748
`define TANH_LUT_NEGATIVE_8750 16'h8750
`define TANH_LUT_NEGATIVE_8758 16'h8758
`define TANH_LUT_NEGATIVE_8760 16'h8760
`define TANH_LUT_NEGATIVE_8768 16'h8768
`define TANH_LUT_NEGATIVE_8770 16'h8770
`define TANH_LUT_NEGATIVE_8778 16'h8778
`define TANH_LUT_NEGATIVE_8780 16'h8780
`define TANH_LUT_NEGATIVE_8788 16'h8788
`define TANH_LUT_NEGATIVE_8790 16'h8790
`define TANH_LUT_NEGATIVE_8798 16'h8798
`define TANH_LUT_NEGATIVE_87A0 16'h87A0
`define TANH_LUT_NEGATIVE_87A8 16'h87A8
`define TANH_LUT_NEGATIVE_87B0 16'h87B0
`define TANH_LUT_NEGATIVE_87B8 16'h87B8
`define TANH_LUT_NEGATIVE_87C0 16'h87C0
`define TANH_LUT_NEGATIVE_87C8 16'h87C8
`define TANH_LUT_NEGATIVE_87D0 16'h87D0
`define TANH_LUT_NEGATIVE_87D8 16'h87D8
`define TANH_LUT_NEGATIVE_87E0 16'h87E0
`define TANH_LUT_NEGATIVE_87E8 16'h87E8
`define TANH_LUT_NEGATIVE_87F0 16'h87F0
`define TANH_LUT_NEGATIVE_87F8 16'h87F8
`define TANH_LUT_NEGATIVE_8800 16'h8800
`define TANH_LUT_NEGATIVE_8808 16'h8808
`define TANH_LUT_NEGATIVE_8810 16'h8810
`define TANH_LUT_NEGATIVE_8818 16'h8818
`define TANH_LUT_NEGATIVE_8820 16'h8820
`define TANH_LUT_NEGATIVE_8828 16'h8828
`define TANH_LUT_NEGATIVE_8830 16'h8830
`define TANH_LUT_NEGATIVE_8838 16'h8838
`define TANH_LUT_NEGATIVE_8840 16'h8840
`define TANH_LUT_NEGATIVE_8848 16'h8848
`define TANH_LUT_NEGATIVE_8850 16'h8850
`define TANH_LUT_NEGATIVE_8858 16'h8858
`define TANH_LUT_NEGATIVE_8860 16'h8860
`define TANH_LUT_NEGATIVE_8868 16'h8868
`define TANH_LUT_NEGATIVE_8870 16'h8870
`define TANH_LUT_NEGATIVE_8878 16'h8878
`define TANH_LUT_NEGATIVE_8880 16'h8880
`define TANH_LUT_NEGATIVE_8888 16'h8888
`define TANH_LUT_NEGATIVE_8890 16'h8890
`define TANH_LUT_NEGATIVE_8898 16'h8898
`define TANH_LUT_NEGATIVE_88A0 16'h88A0
`define TANH_LUT_NEGATIVE_88A8 16'h88A8
`define TANH_LUT_NEGATIVE_88B0 16'h88B0
`define TANH_LUT_NEGATIVE_88B8 16'h88B8
`define TANH_LUT_NEGATIVE_88C0 16'h88C0
`define TANH_LUT_NEGATIVE_88C8 16'h88C8
`define TANH_LUT_NEGATIVE_88D0 16'h88D0
`define TANH_LUT_NEGATIVE_88D8 16'h88D8
`define TANH_LUT_NEGATIVE_88E0 16'h88E0
`define TANH_LUT_NEGATIVE_88E8 16'h88E8
`define TANH_LUT_NEGATIVE_88F0 16'h88F0
`define TANH_LUT_NEGATIVE_88F8 16'h88F8
`define TANH_LUT_NEGATIVE_8900 16'h8900
`define TANH_LUT_NEGATIVE_8908 16'h8908
`define TANH_LUT_NEGATIVE_8910 16'h8910
`define TANH_LUT_NEGATIVE_8918 16'h8918
`define TANH_LUT_NEGATIVE_8920 16'h8920
`define TANH_LUT_NEGATIVE_8928 16'h8928
`define TANH_LUT_NEGATIVE_8930 16'h8930
`define TANH_LUT_NEGATIVE_8938 16'h8938
`define TANH_LUT_NEGATIVE_8940 16'h8940
`define TANH_LUT_NEGATIVE_8948 16'h8948
`define TANH_LUT_NEGATIVE_8950 16'h8950
`define TANH_LUT_NEGATIVE_8958 16'h8958
`define TANH_LUT_NEGATIVE_8960 16'h8960
`define TANH_LUT_NEGATIVE_8968 16'h8968
`define TANH_LUT_NEGATIVE_8970 16'h8970
`define TANH_LUT_NEGATIVE_8978 16'h8978
`define TANH_LUT_NEGATIVE_8980 16'h8980
`define TANH_LUT_NEGATIVE_8988 16'h8988
`define TANH_LUT_NEGATIVE_8990 16'h8990
`define TANH_LUT_NEGATIVE_8998 16'h8998
`define TANH_LUT_NEGATIVE_89A0 16'h89A0
`define TANH_LUT_NEGATIVE_89A8 16'h89A8
`define TANH_LUT_NEGATIVE_89B0 16'h89B0
`define TANH_LUT_NEGATIVE_89B8 16'h89B8
`define TANH_LUT_NEGATIVE_89C0 16'h89C0
`define TANH_LUT_NEGATIVE_89C8 16'h89C8
`define TANH_LUT_NEGATIVE_89D0 16'h89D0
`define TANH_LUT_NEGATIVE_89D8 16'h89D8
`define TANH_LUT_NEGATIVE_89E0 16'h89E0
`define TANH_LUT_NEGATIVE_89E8 16'h89E8
`define TANH_LUT_NEGATIVE_89F0 16'h89F0
`define TANH_LUT_NEGATIVE_89F8 16'h89F8
`define TANH_LUT_NEGATIVE_8A00 16'h8A00
`define TANH_LUT_NEGATIVE_8A08 16'h8A08
`define TANH_LUT_NEGATIVE_8A10 16'h8A10
`define TANH_LUT_NEGATIVE_8A18 16'h8A18
`define TANH_LUT_NEGATIVE_8A20 16'h8A20
`define TANH_LUT_NEGATIVE_8A28 16'h8A28
`define TANH_LUT_NEGATIVE_8A30 16'h8A30
`define TANH_LUT_NEGATIVE_8A38 16'h8A38
`define TANH_LUT_NEGATIVE_8A40 16'h8A40
`define TANH_LUT_NEGATIVE_8A48 16'h8A48
`define TANH_LUT_NEGATIVE_8A50 16'h8A50
`define TANH_LUT_NEGATIVE_8A58 16'h8A58
`define TANH_LUT_NEGATIVE_8A60 16'h8A60
`define TANH_LUT_NEGATIVE_8A68 16'h8A68
`define TANH_LUT_NEGATIVE_8A70 16'h8A70
`define TANH_LUT_NEGATIVE_8A78 16'h8A78
`define TANH_LUT_NEGATIVE_8A80 16'h8A80
`define TANH_LUT_NEGATIVE_8A88 16'h8A88
`define TANH_LUT_NEGATIVE_8A90 16'h8A90
`define TANH_LUT_NEGATIVE_8A98 16'h8A98
`define TANH_LUT_NEGATIVE_8AA0 16'h8AA0
`define TANH_LUT_NEGATIVE_8AA8 16'h8AA8
`define TANH_LUT_NEGATIVE_8AB0 16'h8AB0
`define TANH_LUT_NEGATIVE_8AB8 16'h8AB8
`define TANH_LUT_NEGATIVE_8AC0 16'h8AC0
`define TANH_LUT_NEGATIVE_8AC8 16'h8AC8
`define TANH_LUT_NEGATIVE_8AD0 16'h8AD0
`define TANH_LUT_NEGATIVE_8AD8 16'h8AD8
`define TANH_LUT_NEGATIVE_8AE0 16'h8AE0
`define TANH_LUT_NEGATIVE_8AE8 16'h8AE8
`define TANH_LUT_NEGATIVE_8AF0 16'h8AF0
`define TANH_LUT_NEGATIVE_8AF8 16'h8AF8
`define TANH_LUT_NEGATIVE_8B00 16'h8B00
`define TANH_LUT_NEGATIVE_8B08 16'h8B08
`define TANH_LUT_NEGATIVE_8B10 16'h8B10
`define TANH_LUT_NEGATIVE_8B18 16'h8B18
`define TANH_LUT_NEGATIVE_8B20 16'h8B20
`define TANH_LUT_NEGATIVE_8B28 16'h8B28
`define TANH_LUT_NEGATIVE_8B30 16'h8B30
`define TANH_LUT_NEGATIVE_8B38 16'h8B38
`define TANH_LUT_NEGATIVE_8B40 16'h8B40
`define TANH_LUT_NEGATIVE_8B48 16'h8B48
`define TANH_LUT_NEGATIVE_8B50 16'h8B50
`define TANH_LUT_NEGATIVE_8B58 16'h8B58
`define TANH_LUT_NEGATIVE_8B60 16'h8B60
`define TANH_LUT_NEGATIVE_8B68 16'h8B68
`define TANH_LUT_NEGATIVE_8B70 16'h8B70
`define TANH_LUT_NEGATIVE_8B78 16'h8B78
`define TANH_LUT_NEGATIVE_8B80 16'h8B80
`define TANH_LUT_NEGATIVE_8B88 16'h8B88
`define TANH_LUT_NEGATIVE_8B90 16'h8B90
`define TANH_LUT_NEGATIVE_8B98 16'h8B98
`define TANH_LUT_NEGATIVE_8BA0 16'h8BA0
`define TANH_LUT_NEGATIVE_8BA8 16'h8BA8
`define TANH_LUT_NEGATIVE_8BB0 16'h8BB0
`define TANH_LUT_NEGATIVE_8BB8 16'h8BB8
`define TANH_LUT_NEGATIVE_8BC0 16'h8BC0
`define TANH_LUT_NEGATIVE_8BC8 16'h8BC8
`define TANH_LUT_NEGATIVE_8BD0 16'h8BD0
`define TANH_LUT_NEGATIVE_8BD8 16'h8BD8
`define TANH_LUT_NEGATIVE_8BE0 16'h8BE0
`define TANH_LUT_NEGATIVE_8BE8 16'h8BE8
`define TANH_LUT_NEGATIVE_8BF0 16'h8BF0
`define TANH_LUT_NEGATIVE_8BF8 16'h8BF8
`define TANH_LUT_NEGATIVE_8C00 16'h8C00
`define TANH_LUT_NEGATIVE_8C08 16'h8C08
`define TANH_LUT_NEGATIVE_8C10 16'h8C10
`define TANH_LUT_NEGATIVE_8C18 16'h8C18
`define TANH_LUT_NEGATIVE_8C20 16'h8C20
`define TANH_LUT_NEGATIVE_8C28 16'h8C28
`define TANH_LUT_NEGATIVE_8C30 16'h8C30
`define TANH_LUT_NEGATIVE_8C38 16'h8C38
`define TANH_LUT_NEGATIVE_8C40 16'h8C40
`define TANH_LUT_NEGATIVE_8C48 16'h8C48
`define TANH_LUT_NEGATIVE_8C50 16'h8C50
`define TANH_LUT_NEGATIVE_8C58 16'h8C58
`define TANH_LUT_NEGATIVE_8C60 16'h8C60
`define TANH_LUT_NEGATIVE_8C68 16'h8C68
`define TANH_LUT_NEGATIVE_8C70 16'h8C70
`define TANH_LUT_NEGATIVE_8C78 16'h8C78
`define TANH_LUT_NEGATIVE_8C80 16'h8C80
`define TANH_LUT_NEGATIVE_8C88 16'h8C88
`define TANH_LUT_NEGATIVE_8C90 16'h8C90
`define TANH_LUT_NEGATIVE_8C98 16'h8C98
`define TANH_LUT_NEGATIVE_8CA0 16'h8CA0
`define TANH_LUT_NEGATIVE_8CA8 16'h8CA8
`define TANH_LUT_NEGATIVE_8CB0 16'h8CB0
`define TANH_LUT_NEGATIVE_8CB8 16'h8CB8
`define TANH_LUT_NEGATIVE_8CC0 16'h8CC0
`define TANH_LUT_NEGATIVE_8CC8 16'h8CC8
`define TANH_LUT_NEGATIVE_8CD0 16'h8CD0
`define TANH_LUT_NEGATIVE_8CD8 16'h8CD8
`define TANH_LUT_NEGATIVE_8CE0 16'h8CE0
`define TANH_LUT_NEGATIVE_8CE8 16'h8CE8
`define TANH_LUT_NEGATIVE_8CF0 16'h8CF0
`define TANH_LUT_NEGATIVE_8CF8 16'h8CF8
`define TANH_LUT_NEGATIVE_8D00 16'h8D00
`define TANH_LUT_NEGATIVE_8D08 16'h8D08
`define TANH_LUT_NEGATIVE_8D10 16'h8D10
`define TANH_LUT_NEGATIVE_8D18 16'h8D18
`define TANH_LUT_NEGATIVE_8D20 16'h8D20
`define TANH_LUT_NEGATIVE_8D28 16'h8D28
`define TANH_LUT_NEGATIVE_8D30 16'h8D30
`define TANH_LUT_NEGATIVE_8D38 16'h8D38
`define TANH_LUT_NEGATIVE_8D40 16'h8D40
`define TANH_LUT_NEGATIVE_8D48 16'h8D48
`define TANH_LUT_NEGATIVE_8D50 16'h8D50
`define TANH_LUT_NEGATIVE_8D58 16'h8D58
`define TANH_LUT_NEGATIVE_8D60 16'h8D60
`define TANH_LUT_NEGATIVE_8D68 16'h8D68
`define TANH_LUT_NEGATIVE_8D70 16'h8D70
`define TANH_LUT_NEGATIVE_8D78 16'h8D78
`define TANH_LUT_NEGATIVE_8D80 16'h8D80
`define TANH_LUT_NEGATIVE_8D88 16'h8D88
`define TANH_LUT_NEGATIVE_8D90 16'h8D90
`define TANH_LUT_NEGATIVE_8D98 16'h8D98
`define TANH_LUT_NEGATIVE_8DA0 16'h8DA0
`define TANH_LUT_NEGATIVE_8DA8 16'h8DA8
`define TANH_LUT_NEGATIVE_8DB0 16'h8DB0
`define TANH_LUT_NEGATIVE_8DB8 16'h8DB8
`define TANH_LUT_NEGATIVE_8DC0 16'h8DC0
`define TANH_LUT_NEGATIVE_8DC8 16'h8DC8
`define TANH_LUT_NEGATIVE_8DD0 16'h8DD0
`define TANH_LUT_NEGATIVE_8DD8 16'h8DD8
`define TANH_LUT_NEGATIVE_8DE0 16'h8DE0
`define TANH_LUT_NEGATIVE_8DE8 16'h8DE8
`define TANH_LUT_NEGATIVE_8DF0 16'h8DF0
`define TANH_LUT_NEGATIVE_8DF8 16'h8DF8
`define TANH_LUT_NEGATIVE_8E00 16'h8E00
`define TANH_LUT_NEGATIVE_8E08 16'h8E08
`define TANH_LUT_NEGATIVE_8E10 16'h8E10
`define TANH_LUT_NEGATIVE_8E18 16'h8E18
`define TANH_LUT_NEGATIVE_8E20 16'h8E20
`define TANH_LUT_NEGATIVE_8E28 16'h8E28
`define TANH_LUT_NEGATIVE_8E30 16'h8E30
`define TANH_LUT_NEGATIVE_8E38 16'h8E38
`define TANH_LUT_NEGATIVE_8E40 16'h8E40
`define TANH_LUT_NEGATIVE_8E48 16'h8E48
`define TANH_LUT_NEGATIVE_8E50 16'h8E50
`define TANH_LUT_NEGATIVE_8E58 16'h8E58
`define TANH_LUT_NEGATIVE_8E60 16'h8E60
`define TANH_LUT_NEGATIVE_8E68 16'h8E68
`define TANH_LUT_NEGATIVE_8E70 16'h8E70
`define TANH_LUT_NEGATIVE_8E78 16'h8E78
`define TANH_LUT_NEGATIVE_8E80 16'h8E80
`define TANH_LUT_NEGATIVE_8E88 16'h8E88
`define TANH_LUT_NEGATIVE_8E90 16'h8E90
`define TANH_LUT_NEGATIVE_8E98 16'h8E98
`define TANH_LUT_NEGATIVE_8EA0 16'h8EA0
`define TANH_LUT_NEGATIVE_8EA8 16'h8EA8
`define TANH_LUT_NEGATIVE_8EB0 16'h8EB0
`define TANH_LUT_NEGATIVE_8EB8 16'h8EB8
`define TANH_LUT_NEGATIVE_8EC0 16'h8EC0
`define TANH_LUT_NEGATIVE_8EC8 16'h8EC8
`define TANH_LUT_NEGATIVE_8ED0 16'h8ED0
`define TANH_LUT_NEGATIVE_8ED8 16'h8ED8
`define TANH_LUT_NEGATIVE_8EE0 16'h8EE0
`define TANH_LUT_NEGATIVE_8EE8 16'h8EE8
`define TANH_LUT_NEGATIVE_8EF0 16'h8EF0
`define TANH_LUT_NEGATIVE_8EF8 16'h8EF8
`define TANH_LUT_NEGATIVE_8F00 16'h8F00
`define TANH_LUT_NEGATIVE_8F08 16'h8F08
`define TANH_LUT_NEGATIVE_8F10 16'h8F10
`define TANH_LUT_NEGATIVE_8F18 16'h8F18
`define TANH_LUT_NEGATIVE_8F20 16'h8F20
`define TANH_LUT_NEGATIVE_8F28 16'h8F28
`define TANH_LUT_NEGATIVE_8F30 16'h8F30
`define TANH_LUT_NEGATIVE_8F38 16'h8F38
`define TANH_LUT_NEGATIVE_8F40 16'h8F40
`define TANH_LUT_NEGATIVE_8F48 16'h8F48
`define TANH_LUT_NEGATIVE_8F50 16'h8F50
`define TANH_LUT_NEGATIVE_8F58 16'h8F58
`define TANH_LUT_NEGATIVE_8F60 16'h8F60
`define TANH_LUT_NEGATIVE_8F68 16'h8F68
`define TANH_LUT_NEGATIVE_8F70 16'h8F70
`define TANH_LUT_NEGATIVE_8F78 16'h8F78
`define TANH_LUT_NEGATIVE_8F80 16'h8F80
`define TANH_LUT_NEGATIVE_8F88 16'h8F88
`define TANH_LUT_NEGATIVE_8F90 16'h8F90
`define TANH_LUT_NEGATIVE_8F98 16'h8F98
`define TANH_LUT_NEGATIVE_8FA0 16'h8FA0
`define TANH_LUT_NEGATIVE_8FA8 16'h8FA8
`define TANH_LUT_NEGATIVE_8FB0 16'h8FB0
`define TANH_LUT_NEGATIVE_8FB8 16'h8FB8
`define TANH_LUT_NEGATIVE_8FC0 16'h8FC0
`define TANH_LUT_NEGATIVE_8FC8 16'h8FC8
`define TANH_LUT_NEGATIVE_8FD0 16'h8FD0
`define TANH_LUT_NEGATIVE_8FD8 16'h8FD8
`define TANH_LUT_NEGATIVE_8FE0 16'h8FE0
`define TANH_LUT_NEGATIVE_8FE8 16'h8FE8
`define TANH_LUT_NEGATIVE_8FF0 16'h8FF0
`define TANH_LUT_NEGATIVE_8FF8 16'h8FF8
`define TANH_LUT_NEGATIVE_9000 16'h9000
`define TANH_LUT_NEGATIVE_9008 16'h9008
`define TANH_LUT_NEGATIVE_9010 16'h9010
`define TANH_LUT_NEGATIVE_9018 16'h9018
`define TANH_LUT_NEGATIVE_9020 16'h9020
`define TANH_LUT_NEGATIVE_9028 16'h9028
`define TANH_LUT_NEGATIVE_9030 16'h9030
`define TANH_LUT_NEGATIVE_9038 16'h9038
`define TANH_LUT_NEGATIVE_9040 16'h9040
`define TANH_LUT_NEGATIVE_9048 16'h9048
`define TANH_LUT_NEGATIVE_9050 16'h9050
`define TANH_LUT_NEGATIVE_9058 16'h9058
`define TANH_LUT_NEGATIVE_9060 16'h9060
`define TANH_LUT_NEGATIVE_9068 16'h9068
`define TANH_LUT_NEGATIVE_9070 16'h9070
`define TANH_LUT_NEGATIVE_9078 16'h9078
`define TANH_LUT_NEGATIVE_9080 16'h9080
`define TANH_LUT_NEGATIVE_9088 16'h9088
`define TANH_LUT_NEGATIVE_9090 16'h9090
`define TANH_LUT_NEGATIVE_9098 16'h9098
`define TANH_LUT_NEGATIVE_90A0 16'h90A0
`define TANH_LUT_NEGATIVE_90A8 16'h90A8
`define TANH_LUT_NEGATIVE_90B0 16'h90B0
`define TANH_LUT_NEGATIVE_90B8 16'h90B8
`define TANH_LUT_NEGATIVE_90C0 16'h90C0
`define TANH_LUT_NEGATIVE_90C8 16'h90C8
`define TANH_LUT_NEGATIVE_90D0 16'h90D0
`define TANH_LUT_NEGATIVE_90D8 16'h90D8
`define TANH_LUT_NEGATIVE_90E0 16'h90E0
`define TANH_LUT_NEGATIVE_90E8 16'h90E8
`define TANH_LUT_NEGATIVE_90F0 16'h90F0
`define TANH_LUT_NEGATIVE_90F8 16'h90F8
`define TANH_LUT_NEGATIVE_9100 16'h9100
`define TANH_LUT_NEGATIVE_9108 16'h9108
`define TANH_LUT_NEGATIVE_9110 16'h9110
`define TANH_LUT_NEGATIVE_9118 16'h9118
`define TANH_LUT_NEGATIVE_9120 16'h9120
`define TANH_LUT_NEGATIVE_9128 16'h9128
`define TANH_LUT_NEGATIVE_9130 16'h9130
`define TANH_LUT_NEGATIVE_9138 16'h9138
`define TANH_LUT_NEGATIVE_9140 16'h9140
`define TANH_LUT_NEGATIVE_9148 16'h9148
`define TANH_LUT_NEGATIVE_9150 16'h9150
`define TANH_LUT_NEGATIVE_9158 16'h9158
`define TANH_LUT_NEGATIVE_9160 16'h9160
`define TANH_LUT_NEGATIVE_9168 16'h9168
`define TANH_LUT_NEGATIVE_9170 16'h9170
`define TANH_LUT_NEGATIVE_9178 16'h9178
`define TANH_LUT_NEGATIVE_9180 16'h9180
`define TANH_LUT_NEGATIVE_9188 16'h9188
`define TANH_LUT_NEGATIVE_9190 16'h9190
`define TANH_LUT_NEGATIVE_9198 16'h9198
`define TANH_LUT_NEGATIVE_91A0 16'h91A0
`define TANH_LUT_NEGATIVE_91A8 16'h91A8
`define TANH_LUT_NEGATIVE_91B0 16'h91B0
`define TANH_LUT_NEGATIVE_91B8 16'h91B8
`define TANH_LUT_NEGATIVE_91C0 16'h91C0
`define TANH_LUT_NEGATIVE_91C8 16'h91C8
`define TANH_LUT_NEGATIVE_91D0 16'h91D0
`define TANH_LUT_NEGATIVE_91D8 16'h91D8
`define TANH_LUT_NEGATIVE_91E0 16'h91E0
`define TANH_LUT_NEGATIVE_91E8 16'h91E8
`define TANH_LUT_NEGATIVE_91F0 16'h91F0
`define TANH_LUT_NEGATIVE_91F8 16'h91F8
`define TANH_LUT_NEGATIVE_9200 16'h9200
`define TANH_LUT_NEGATIVE_9208 16'h9208
`define TANH_LUT_NEGATIVE_9210 16'h9210
`define TANH_LUT_NEGATIVE_9218 16'h9218
`define TANH_LUT_NEGATIVE_9220 16'h9220
`define TANH_LUT_NEGATIVE_9228 16'h9228
`define TANH_LUT_NEGATIVE_9230 16'h9230
`define TANH_LUT_NEGATIVE_9238 16'h9238
`define TANH_LUT_NEGATIVE_9240 16'h9240
`define TANH_LUT_NEGATIVE_9248 16'h9248
`define TANH_LUT_NEGATIVE_9250 16'h9250
`define TANH_LUT_NEGATIVE_9258 16'h9258
`define TANH_LUT_NEGATIVE_9260 16'h9260
`define TANH_LUT_NEGATIVE_9268 16'h9268
`define TANH_LUT_NEGATIVE_9270 16'h9270
`define TANH_LUT_NEGATIVE_9278 16'h9278
`define TANH_LUT_NEGATIVE_9280 16'h9280
`define TANH_LUT_NEGATIVE_9288 16'h9288
`define TANH_LUT_NEGATIVE_9290 16'h9290
`define TANH_LUT_NEGATIVE_9298 16'h9298
`define TANH_LUT_NEGATIVE_92A0 16'h92A0
`define TANH_LUT_NEGATIVE_92A8 16'h92A8
`define TANH_LUT_NEGATIVE_92B0 16'h92B0
`define TANH_LUT_NEGATIVE_92B8 16'h92B8
`define TANH_LUT_NEGATIVE_92C0 16'h92C0
`define TANH_LUT_NEGATIVE_92C8 16'h92C8
`define TANH_LUT_NEGATIVE_92D0 16'h92D0
`define TANH_LUT_NEGATIVE_92D8 16'h92D8
`define TANH_LUT_NEGATIVE_92E0 16'h92E0
`define TANH_LUT_NEGATIVE_92E8 16'h92E8
`define TANH_LUT_NEGATIVE_92F0 16'h92F0
`define TANH_LUT_NEGATIVE_92F8 16'h92F8
`define TANH_LUT_NEGATIVE_9300 16'h9300
`define TANH_LUT_NEGATIVE_9308 16'h9308
`define TANH_LUT_NEGATIVE_9310 16'h9310
`define TANH_LUT_NEGATIVE_9318 16'h9318
`define TANH_LUT_NEGATIVE_9320 16'h9320
`define TANH_LUT_NEGATIVE_9328 16'h9328
`define TANH_LUT_NEGATIVE_9330 16'h9330
`define TANH_LUT_NEGATIVE_9338 16'h9338
`define TANH_LUT_NEGATIVE_9340 16'h9340
`define TANH_LUT_NEGATIVE_9348 16'h9348
`define TANH_LUT_NEGATIVE_9350 16'h9350
`define TANH_LUT_NEGATIVE_9358 16'h9358
`define TANH_LUT_NEGATIVE_9360 16'h9360
`define TANH_LUT_NEGATIVE_9368 16'h9368
`define TANH_LUT_NEGATIVE_9370 16'h9370
`define TANH_LUT_NEGATIVE_9378 16'h9378
`define TANH_LUT_NEGATIVE_9380 16'h9380
`define TANH_LUT_NEGATIVE_9388 16'h9388
`define TANH_LUT_NEGATIVE_9390 16'h9390
`define TANH_LUT_NEGATIVE_9398 16'h9398
`define TANH_LUT_NEGATIVE_93A0 16'h93A0
`define TANH_LUT_NEGATIVE_93A8 16'h93A8
`define TANH_LUT_NEGATIVE_93B0 16'h93B0
`define TANH_LUT_NEGATIVE_93B8 16'h93B8
`define TANH_LUT_NEGATIVE_93C0 16'h93C0
`define TANH_LUT_NEGATIVE_93C8 16'h93C8
`define TANH_LUT_NEGATIVE_93D0 16'h93D0
`define TANH_LUT_NEGATIVE_93D8 16'h93D8
`define TANH_LUT_NEGATIVE_93E0 16'h93E0
`define TANH_LUT_NEGATIVE_93E8 16'h93E8
`define TANH_LUT_NEGATIVE_93F0 16'h93F0
`define TANH_LUT_NEGATIVE_93F8 16'h93F8
`define TANH_LUT_NEGATIVE_9400 16'h9400
`define TANH_LUT_NEGATIVE_9408 16'h9408
`define TANH_LUT_NEGATIVE_9410 16'h9410
`define TANH_LUT_NEGATIVE_9418 16'h9418
`define TANH_LUT_NEGATIVE_9420 16'h9420
`define TANH_LUT_NEGATIVE_9428 16'h9428
`define TANH_LUT_NEGATIVE_9430 16'h9430
`define TANH_LUT_NEGATIVE_9438 16'h9438
`define TANH_LUT_NEGATIVE_9440 16'h9440
`define TANH_LUT_NEGATIVE_9448 16'h9448
`define TANH_LUT_NEGATIVE_9450 16'h9450
`define TANH_LUT_NEGATIVE_9458 16'h9458
`define TANH_LUT_NEGATIVE_9460 16'h9460
`define TANH_LUT_NEGATIVE_9468 16'h9468
`define TANH_LUT_NEGATIVE_9470 16'h9470
`define TANH_LUT_NEGATIVE_9478 16'h9478
`define TANH_LUT_NEGATIVE_9480 16'h9480
`define TANH_LUT_NEGATIVE_9488 16'h9488
`define TANH_LUT_NEGATIVE_9490 16'h9490
`define TANH_LUT_NEGATIVE_9498 16'h9498
`define TANH_LUT_NEGATIVE_94A0 16'h94A0
`define TANH_LUT_NEGATIVE_94A8 16'h94A8
`define TANH_LUT_NEGATIVE_94B0 16'h94B0
`define TANH_LUT_NEGATIVE_94B8 16'h94B8
`define TANH_LUT_NEGATIVE_94C0 16'h94C0
`define TANH_LUT_NEGATIVE_94C8 16'h94C8
`define TANH_LUT_NEGATIVE_94D0 16'h94D0
`define TANH_LUT_NEGATIVE_94D8 16'h94D8
`define TANH_LUT_NEGATIVE_94E0 16'h94E0
`define TANH_LUT_NEGATIVE_94E8 16'h94E8
`define TANH_LUT_NEGATIVE_94F0 16'h94F0
`define TANH_LUT_NEGATIVE_94F8 16'h94F8
`define TANH_LUT_NEGATIVE_9500 16'h9500
`define TANH_LUT_NEGATIVE_9508 16'h9508
`define TANH_LUT_NEGATIVE_9510 16'h9510
`define TANH_LUT_NEGATIVE_9518 16'h9518
`define TANH_LUT_NEGATIVE_9520 16'h9520
`define TANH_LUT_NEGATIVE_9528 16'h9528
`define TANH_LUT_NEGATIVE_9530 16'h9530
`define TANH_LUT_NEGATIVE_9538 16'h9538
`define TANH_LUT_NEGATIVE_9540 16'h9540
`define TANH_LUT_NEGATIVE_9548 16'h9548
`define TANH_LUT_NEGATIVE_9550 16'h9550
`define TANH_LUT_NEGATIVE_9558 16'h9558
`define TANH_LUT_NEGATIVE_9560 16'h9560
`define TANH_LUT_NEGATIVE_9568 16'h9568
`define TANH_LUT_NEGATIVE_9570 16'h9570
`define TANH_LUT_NEGATIVE_9578 16'h9578
`define TANH_LUT_NEGATIVE_9580 16'h9580
`define TANH_LUT_NEGATIVE_9588 16'h9588
`define TANH_LUT_NEGATIVE_9590 16'h9590
`define TANH_LUT_NEGATIVE_9598 16'h9598
`define TANH_LUT_NEGATIVE_95A0 16'h95A0
`define TANH_LUT_NEGATIVE_95A8 16'h95A8
`define TANH_LUT_NEGATIVE_95B0 16'h95B0
`define TANH_LUT_NEGATIVE_95B8 16'h95B8
`define TANH_LUT_NEGATIVE_95C0 16'h95C0
`define TANH_LUT_NEGATIVE_95C8 16'h95C8
`define TANH_LUT_NEGATIVE_95D0 16'h95D0
`define TANH_LUT_NEGATIVE_95D8 16'h95D8
`define TANH_LUT_NEGATIVE_95E0 16'h95E0
`define TANH_LUT_NEGATIVE_95E8 16'h95E8
`define TANH_LUT_NEGATIVE_95F0 16'h95F0
`define TANH_LUT_NEGATIVE_95F8 16'h95F8
`define TANH_LUT_NEGATIVE_9600 16'h9600
`define TANH_LUT_NEGATIVE_9608 16'h9608
`define TANH_LUT_NEGATIVE_9610 16'h9610
`define TANH_LUT_NEGATIVE_9618 16'h9618
`define TANH_LUT_NEGATIVE_9620 16'h9620
`define TANH_LUT_NEGATIVE_9628 16'h9628
`define TANH_LUT_NEGATIVE_9630 16'h9630
`define TANH_LUT_NEGATIVE_9638 16'h9638
`define TANH_LUT_NEGATIVE_9640 16'h9640
`define TANH_LUT_NEGATIVE_9648 16'h9648
`define TANH_LUT_NEGATIVE_9650 16'h9650
`define TANH_LUT_NEGATIVE_9658 16'h9658
`define TANH_LUT_NEGATIVE_9660 16'h9660
`define TANH_LUT_NEGATIVE_9668 16'h9668
`define TANH_LUT_NEGATIVE_9670 16'h9670
`define TANH_LUT_NEGATIVE_9678 16'h9678
`define TANH_LUT_NEGATIVE_9680 16'h9680
`define TANH_LUT_NEGATIVE_9688 16'h9688
`define TANH_LUT_NEGATIVE_9690 16'h9690
`define TANH_LUT_NEGATIVE_9698 16'h9698
`define TANH_LUT_NEGATIVE_96A0 16'h96A0
`define TANH_LUT_NEGATIVE_96A8 16'h96A8
`define TANH_LUT_NEGATIVE_96B0 16'h96B0
`define TANH_LUT_NEGATIVE_96B8 16'h96B8
`define TANH_LUT_NEGATIVE_96C0 16'h96C0
`define TANH_LUT_NEGATIVE_96C8 16'h96C8
`define TANH_LUT_NEGATIVE_96D0 16'h96D0
`define TANH_LUT_NEGATIVE_96D8 16'h96D8
`define TANH_LUT_NEGATIVE_96E0 16'h96E0
`define TANH_LUT_NEGATIVE_96E8 16'h96E8
`define TANH_LUT_NEGATIVE_96F0 16'h96F0
`define TANH_LUT_NEGATIVE_96F8 16'h96F8
`define TANH_LUT_NEGATIVE_9700 16'h9700
`define TANH_LUT_NEGATIVE_9708 16'h9708
`define TANH_LUT_NEGATIVE_9710 16'h9710
`define TANH_LUT_NEGATIVE_9718 16'h9718
`define TANH_LUT_NEGATIVE_9720 16'h9720
`define TANH_LUT_NEGATIVE_9728 16'h9728
`define TANH_LUT_NEGATIVE_9730 16'h9730
`define TANH_LUT_NEGATIVE_9738 16'h9738
`define TANH_LUT_NEGATIVE_9740 16'h9740
`define TANH_LUT_NEGATIVE_9748 16'h9748
`define TANH_LUT_NEGATIVE_9750 16'h9750
`define TANH_LUT_NEGATIVE_9758 16'h9758
`define TANH_LUT_NEGATIVE_9760 16'h9760
`define TANH_LUT_NEGATIVE_9768 16'h9768
`define TANH_LUT_NEGATIVE_9770 16'h9770
`define TANH_LUT_NEGATIVE_9778 16'h9778
`define TANH_LUT_NEGATIVE_9780 16'h9780
`define TANH_LUT_NEGATIVE_9788 16'h9788
`define TANH_LUT_NEGATIVE_9790 16'h9790
`define TANH_LUT_NEGATIVE_9798 16'h9798
`define TANH_LUT_NEGATIVE_97A0 16'h97A0
`define TANH_LUT_NEGATIVE_97A8 16'h97A8
`define TANH_LUT_NEGATIVE_97B0 16'h97B0
`define TANH_LUT_NEGATIVE_97B8 16'h97B8
`define TANH_LUT_NEGATIVE_97C0 16'h97C0
`define TANH_LUT_NEGATIVE_97C8 16'h97C8
`define TANH_LUT_NEGATIVE_97D0 16'h97D0
`define TANH_LUT_NEGATIVE_97D8 16'h97D8
`define TANH_LUT_NEGATIVE_97E0 16'h97E0
`define TANH_LUT_NEGATIVE_97E8 16'h97E8
`define TANH_LUT_NEGATIVE_97F0 16'h97F0
`define TANH_LUT_NEGATIVE_97F8 16'h97F8
`define TANH_LUT_NEGATIVE_9800 16'h9800
`define TANH_LUT_NEGATIVE_9808 16'h9808
`define TANH_LUT_NEGATIVE_9810 16'h9810
`define TANH_LUT_NEGATIVE_9818 16'h9818
`define TANH_LUT_NEGATIVE_9820 16'h9820
`define TANH_LUT_NEGATIVE_9828 16'h9828
`define TANH_LUT_NEGATIVE_9830 16'h9830
`define TANH_LUT_NEGATIVE_9838 16'h9838
`define TANH_LUT_NEGATIVE_9840 16'h9840
`define TANH_LUT_NEGATIVE_9848 16'h9848
`define TANH_LUT_NEGATIVE_9850 16'h9850
`define TANH_LUT_NEGATIVE_9858 16'h9858
`define TANH_LUT_NEGATIVE_9860 16'h9860
`define TANH_LUT_NEGATIVE_9868 16'h9868
`define TANH_LUT_NEGATIVE_9870 16'h9870
`define TANH_LUT_NEGATIVE_9878 16'h9878
`define TANH_LUT_NEGATIVE_9880 16'h9880
`define TANH_LUT_NEGATIVE_9888 16'h9888
`define TANH_LUT_NEGATIVE_9890 16'h9890
`define TANH_LUT_NEGATIVE_9898 16'h9898
`define TANH_LUT_NEGATIVE_98A0 16'h98A0
`define TANH_LUT_NEGATIVE_98A8 16'h98A8
`define TANH_LUT_NEGATIVE_98B0 16'h98B0
`define TANH_LUT_NEGATIVE_98B8 16'h98B8
`define TANH_LUT_NEGATIVE_98C0 16'h98C0
`define TANH_LUT_NEGATIVE_98C8 16'h98C8
`define TANH_LUT_NEGATIVE_98D0 16'h98D0
`define TANH_LUT_NEGATIVE_98D8 16'h98D8
`define TANH_LUT_NEGATIVE_98E0 16'h98E0
`define TANH_LUT_NEGATIVE_98E8 16'h98E8
`define TANH_LUT_NEGATIVE_98F0 16'h98F0
`define TANH_LUT_NEGATIVE_98F8 16'h98F8
`define TANH_LUT_NEGATIVE_9900 16'h9900
`define TANH_LUT_NEGATIVE_9908 16'h9908
`define TANH_LUT_NEGATIVE_9910 16'h9910
`define TANH_LUT_NEGATIVE_9918 16'h9918
`define TANH_LUT_NEGATIVE_9920 16'h9920
`define TANH_LUT_NEGATIVE_9928 16'h9928
`define TANH_LUT_NEGATIVE_9930 16'h9930
`define TANH_LUT_NEGATIVE_9938 16'h9938
`define TANH_LUT_NEGATIVE_9940 16'h9940
`define TANH_LUT_NEGATIVE_9948 16'h9948
`define TANH_LUT_NEGATIVE_9950 16'h9950
`define TANH_LUT_NEGATIVE_9958 16'h9958
`define TANH_LUT_NEGATIVE_9960 16'h9960
`define TANH_LUT_NEGATIVE_9968 16'h9968
`define TANH_LUT_NEGATIVE_9970 16'h9970
`define TANH_LUT_NEGATIVE_9978 16'h9978
`define TANH_LUT_NEGATIVE_9980 16'h9980
`define TANH_LUT_NEGATIVE_9988 16'h9988
`define TANH_LUT_NEGATIVE_9990 16'h9990
`define TANH_LUT_NEGATIVE_9998 16'h9998
`define TANH_LUT_NEGATIVE_99A0 16'h99A0
`define TANH_LUT_NEGATIVE_99A8 16'h99A8
`define TANH_LUT_NEGATIVE_99B0 16'h99B0
`define TANH_LUT_NEGATIVE_99B8 16'h99B8
`define TANH_LUT_NEGATIVE_99C0 16'h99C0
`define TANH_LUT_NEGATIVE_99C8 16'h99C8
`define TANH_LUT_NEGATIVE_99D0 16'h99D0
`define TANH_LUT_NEGATIVE_99D8 16'h99D8
`define TANH_LUT_NEGATIVE_99E0 16'h99E0
`define TANH_LUT_NEGATIVE_99E8 16'h99E8
`define TANH_LUT_NEGATIVE_99F0 16'h99F0
`define TANH_LUT_NEGATIVE_99F8 16'h99F8
`define TANH_LUT_NEGATIVE_9A00 16'h9A00
`define TANH_LUT_NEGATIVE_9A08 16'h9A08
`define TANH_LUT_NEGATIVE_9A10 16'h9A10
`define TANH_LUT_NEGATIVE_9A18 16'h9A18
`define TANH_LUT_NEGATIVE_9A20 16'h9A20
`define TANH_LUT_NEGATIVE_9A28 16'h9A28
`define TANH_LUT_NEGATIVE_9A30 16'h9A30
`define TANH_LUT_NEGATIVE_9A38 16'h9A38
`define TANH_LUT_NEGATIVE_9A40 16'h9A40
`define TANH_LUT_NEGATIVE_9A48 16'h9A48
`define TANH_LUT_NEGATIVE_9A50 16'h9A50
`define TANH_LUT_NEGATIVE_9A58 16'h9A58
`define TANH_LUT_NEGATIVE_9A60 16'h9A60
`define TANH_LUT_NEGATIVE_9A68 16'h9A68
`define TANH_LUT_NEGATIVE_9A70 16'h9A70
`define TANH_LUT_NEGATIVE_9A78 16'h9A78
`define TANH_LUT_NEGATIVE_9A80 16'h9A80
`define TANH_LUT_NEGATIVE_9A88 16'h9A88
`define TANH_LUT_NEGATIVE_9A90 16'h9A90
`define TANH_LUT_NEGATIVE_9A98 16'h9A98
`define TANH_LUT_NEGATIVE_9AA0 16'h9AA0
`define TANH_LUT_NEGATIVE_9AA8 16'h9AA8
`define TANH_LUT_NEGATIVE_9AB0 16'h9AB0
`define TANH_LUT_NEGATIVE_9AB8 16'h9AB8
`define TANH_LUT_NEGATIVE_9AC0 16'h9AC0
`define TANH_LUT_NEGATIVE_9AC8 16'h9AC8
`define TANH_LUT_NEGATIVE_9AD0 16'h9AD0
`define TANH_LUT_NEGATIVE_9AD8 16'h9AD8
`define TANH_LUT_NEGATIVE_9AE0 16'h9AE0
`define TANH_LUT_NEGATIVE_9AE8 16'h9AE8
`define TANH_LUT_NEGATIVE_9AF0 16'h9AF0
`define TANH_LUT_NEGATIVE_9AF8 16'h9AF8
`define TANH_LUT_NEGATIVE_9B00 16'h9B00
`define TANH_LUT_NEGATIVE_9B08 16'h9B08
`define TANH_LUT_NEGATIVE_9B10 16'h9B10
`define TANH_LUT_NEGATIVE_9B18 16'h9B18
`define TANH_LUT_NEGATIVE_9B20 16'h9B20
`define TANH_LUT_NEGATIVE_9B28 16'h9B28
`define TANH_LUT_NEGATIVE_9B30 16'h9B30
`define TANH_LUT_NEGATIVE_9B38 16'h9B38
`define TANH_LUT_NEGATIVE_9B40 16'h9B40
`define TANH_LUT_NEGATIVE_9B48 16'h9B48
`define TANH_LUT_NEGATIVE_9B50 16'h9B50
`define TANH_LUT_NEGATIVE_9B58 16'h9B58
`define TANH_LUT_NEGATIVE_9B60 16'h9B60
`define TANH_LUT_NEGATIVE_9B68 16'h9B68
`define TANH_LUT_NEGATIVE_9B70 16'h9B70
`define TANH_LUT_NEGATIVE_9B78 16'h9B78
`define TANH_LUT_NEGATIVE_9B80 16'h9B80
`define TANH_LUT_NEGATIVE_9B88 16'h9B88
`define TANH_LUT_NEGATIVE_9B90 16'h9B90
`define TANH_LUT_NEGATIVE_9B98 16'h9B98
`define TANH_LUT_NEGATIVE_9BA0 16'h9BA0
`define TANH_LUT_NEGATIVE_9BA8 16'h9BA8
`define TANH_LUT_NEGATIVE_9BB0 16'h9BB0
`define TANH_LUT_NEGATIVE_9BB8 16'h9BB8
`define TANH_LUT_NEGATIVE_9BC0 16'h9BC0
`define TANH_LUT_NEGATIVE_9BC8 16'h9BC8
`define TANH_LUT_NEGATIVE_9BD0 16'h9BD0
`define TANH_LUT_NEGATIVE_9BD8 16'h9BD8
`define TANH_LUT_NEGATIVE_9BE0 16'h9BE0
`define TANH_LUT_NEGATIVE_9BE8 16'h9BE8
`define TANH_LUT_NEGATIVE_9BF0 16'h9BF0
`define TANH_LUT_NEGATIVE_9BF8 16'h9BF8
`define TANH_LUT_NEGATIVE_9C00 16'h9C00
`define TANH_LUT_NEGATIVE_9C08 16'h9C08
`define TANH_LUT_NEGATIVE_9C10 16'h9C10
`define TANH_LUT_NEGATIVE_9C18 16'h9C18
`define TANH_LUT_NEGATIVE_9C20 16'h9C20
`define TANH_LUT_NEGATIVE_9C28 16'h9C28
`define TANH_LUT_NEGATIVE_9C30 16'h9C30
`define TANH_LUT_NEGATIVE_9C38 16'h9C38
`define TANH_LUT_NEGATIVE_9C40 16'h9C40
`define TANH_LUT_NEGATIVE_9C48 16'h9C48
`define TANH_LUT_NEGATIVE_9C50 16'h9C50
`define TANH_LUT_NEGATIVE_9C58 16'h9C58
`define TANH_LUT_NEGATIVE_9C60 16'h9C60
`define TANH_LUT_NEGATIVE_9C68 16'h9C68
`define TANH_LUT_NEGATIVE_9C70 16'h9C70
`define TANH_LUT_NEGATIVE_9C78 16'h9C78
`define TANH_LUT_NEGATIVE_9C80 16'h9C80
`define TANH_LUT_NEGATIVE_9C88 16'h9C88
`define TANH_LUT_NEGATIVE_9C90 16'h9C90
`define TANH_LUT_NEGATIVE_9C98 16'h9C98
`define TANH_LUT_NEGATIVE_9CA0 16'h9CA0
`define TANH_LUT_NEGATIVE_9CA8 16'h9CA8
`define TANH_LUT_NEGATIVE_9CB0 16'h9CB0
`define TANH_LUT_NEGATIVE_9CB8 16'h9CB8
`define TANH_LUT_NEGATIVE_9CC0 16'h9CC0
`define TANH_LUT_NEGATIVE_9CC8 16'h9CC8
`define TANH_LUT_NEGATIVE_9CD0 16'h9CD0
`define TANH_LUT_NEGATIVE_9CD8 16'h9CD8
`define TANH_LUT_NEGATIVE_9CE0 16'h9CE0
`define TANH_LUT_NEGATIVE_9CE8 16'h9CE8
`define TANH_LUT_NEGATIVE_9CF0 16'h9CF0
`define TANH_LUT_NEGATIVE_9CF8 16'h9CF8
`define TANH_LUT_NEGATIVE_9D00 16'h9D00
`define TANH_LUT_NEGATIVE_9D08 16'h9D08
`define TANH_LUT_NEGATIVE_9D10 16'h9D10
`define TANH_LUT_NEGATIVE_9D18 16'h9D18
`define TANH_LUT_NEGATIVE_9D20 16'h9D20
`define TANH_LUT_NEGATIVE_9D28 16'h9D28
`define TANH_LUT_NEGATIVE_9D30 16'h9D30
`define TANH_LUT_NEGATIVE_9D38 16'h9D38
`define TANH_LUT_NEGATIVE_9D40 16'h9D40
`define TANH_LUT_NEGATIVE_9D48 16'h9D48
`define TANH_LUT_NEGATIVE_9D50 16'h9D50
`define TANH_LUT_NEGATIVE_9D58 16'h9D58
`define TANH_LUT_NEGATIVE_9D60 16'h9D60
`define TANH_LUT_NEGATIVE_9D68 16'h9D68
`define TANH_LUT_NEGATIVE_9D70 16'h9D70
`define TANH_LUT_NEGATIVE_9D78 16'h9D78
`define TANH_LUT_NEGATIVE_9D80 16'h9D80
`define TANH_LUT_NEGATIVE_9D88 16'h9D88
`define TANH_LUT_NEGATIVE_9D90 16'h9D90
`define TANH_LUT_NEGATIVE_9D98 16'h9D98
`define TANH_LUT_NEGATIVE_9DA0 16'h9DA0
`define TANH_LUT_NEGATIVE_9DA8 16'h9DA8
`define TANH_LUT_NEGATIVE_9DB0 16'h9DB0
`define TANH_LUT_NEGATIVE_9DB8 16'h9DB8
`define TANH_LUT_NEGATIVE_9DC0 16'h9DC0
`define TANH_LUT_NEGATIVE_9DC8 16'h9DC8
`define TANH_LUT_NEGATIVE_9DD0 16'h9DD0
`define TANH_LUT_NEGATIVE_9DD8 16'h9DD8
`define TANH_LUT_NEGATIVE_9DE0 16'h9DE0
`define TANH_LUT_NEGATIVE_9DE8 16'h9DE8
`define TANH_LUT_NEGATIVE_9DF0 16'h9DF0
`define TANH_LUT_NEGATIVE_9DF8 16'h9DF8
`define TANH_LUT_NEGATIVE_9E00 16'h9E00
`define TANH_LUT_NEGATIVE_9E08 16'h9E08
`define TANH_LUT_NEGATIVE_9E10 16'h9E10
`define TANH_LUT_NEGATIVE_9E18 16'h9E18
`define TANH_LUT_NEGATIVE_9E20 16'h9E20
`define TANH_LUT_NEGATIVE_9E28 16'h9E28
`define TANH_LUT_NEGATIVE_9E30 16'h9E30
`define TANH_LUT_NEGATIVE_9E38 16'h9E38
`define TANH_LUT_NEGATIVE_9E40 16'h9E40
`define TANH_LUT_NEGATIVE_9E48 16'h9E48
`define TANH_LUT_NEGATIVE_9E50 16'h9E50
`define TANH_LUT_NEGATIVE_9E58 16'h9E58
`define TANH_LUT_NEGATIVE_9E60 16'h9E60
`define TANH_LUT_NEGATIVE_9E68 16'h9E68
`define TANH_LUT_NEGATIVE_9E70 16'h9E70
`define TANH_LUT_NEGATIVE_9E78 16'h9E78
`define TANH_LUT_NEGATIVE_9E80 16'h9E80
`define TANH_LUT_NEGATIVE_9E88 16'h9E88
`define TANH_LUT_NEGATIVE_9E90 16'h9E90
`define TANH_LUT_NEGATIVE_9E98 16'h9E98
`define TANH_LUT_NEGATIVE_9EA0 16'h9EA0
`define TANH_LUT_NEGATIVE_9EA8 16'h9EA8
`define TANH_LUT_NEGATIVE_9EB0 16'h9EB0
`define TANH_LUT_NEGATIVE_9EB8 16'h9EB8
`define TANH_LUT_NEGATIVE_9EC0 16'h9EC0
`define TANH_LUT_NEGATIVE_9EC8 16'h9EC8
`define TANH_LUT_NEGATIVE_9ED0 16'h9ED0
`define TANH_LUT_NEGATIVE_9ED8 16'h9ED8
`define TANH_LUT_NEGATIVE_9EE0 16'h9EE0
`define TANH_LUT_NEGATIVE_9EE8 16'h9EE8
`define TANH_LUT_NEGATIVE_9EF0 16'h9EF0
`define TANH_LUT_NEGATIVE_9EF8 16'h9EF8
`define TANH_LUT_NEGATIVE_9F00 16'h9F00
`define TANH_LUT_NEGATIVE_9F08 16'h9F08
`define TANH_LUT_NEGATIVE_9F10 16'h9F10
`define TANH_LUT_NEGATIVE_9F18 16'h9F18
`define TANH_LUT_NEGATIVE_9F20 16'h9F20
`define TANH_LUT_NEGATIVE_9F28 16'h9F28
`define TANH_LUT_NEGATIVE_9F30 16'h9F30
`define TANH_LUT_NEGATIVE_9F38 16'h9F38
`define TANH_LUT_NEGATIVE_9F40 16'h9F40
`define TANH_LUT_NEGATIVE_9F48 16'h9F48
`define TANH_LUT_NEGATIVE_9F50 16'h9F50
`define TANH_LUT_NEGATIVE_9F58 16'h9F58
`define TANH_LUT_NEGATIVE_9F60 16'h9F60
`define TANH_LUT_NEGATIVE_9F68 16'h9F68
`define TANH_LUT_NEGATIVE_9F70 16'h9F70
`define TANH_LUT_NEGATIVE_9F78 16'h9F78
`define TANH_LUT_NEGATIVE_9F80 16'h9F80
`define TANH_LUT_NEGATIVE_9F88 16'h9F88
`define TANH_LUT_NEGATIVE_9F90 16'h9F90
`define TANH_LUT_NEGATIVE_9F98 16'h9F98
`define TANH_LUT_NEGATIVE_9FA0 16'h9FA0
`define TANH_LUT_NEGATIVE_9FA8 16'h9FA8
`define TANH_LUT_NEGATIVE_9FB0 16'h9FB0
`define TANH_LUT_NEGATIVE_9FB8 16'h9FB8
`define TANH_LUT_NEGATIVE_9FC0 16'h9FC0
`define TANH_LUT_NEGATIVE_9FC8 16'h9FC8
`define TANH_LUT_NEGATIVE_9FD0 16'h9FD0
`define TANH_LUT_NEGATIVE_9FD8 16'h9FD8
`define TANH_LUT_NEGATIVE_9FE0 16'h9FE0
`define TANH_LUT_NEGATIVE_9FE8 16'h9FE8
`define TANH_LUT_NEGATIVE_9FF0 16'h9FF0
`define TANH_LUT_NEGATIVE_9FF8 16'h9FF8
`define TANH_LUT_NEGATIVE_A000 16'hA000
`define TANH_LUT_NEGATIVE_A008 16'hA008
`define TANH_LUT_NEGATIVE_A010 16'hA010
`define TANH_LUT_NEGATIVE_A018 16'hA018
`define TANH_LUT_NEGATIVE_A020 16'hA020
`define TANH_LUT_NEGATIVE_A028 16'hA028
`define TANH_LUT_NEGATIVE_A030 16'hA030
`define TANH_LUT_NEGATIVE_A038 16'hA038
`define TANH_LUT_NEGATIVE_A040 16'hA040
`define TANH_LUT_NEGATIVE_A048 16'hA048
`define TANH_LUT_NEGATIVE_A050 16'hA050
`define TANH_LUT_NEGATIVE_A058 16'hA058
`define TANH_LUT_NEGATIVE_A060 16'hA060
`define TANH_LUT_NEGATIVE_A068 16'hA068
`define TANH_LUT_NEGATIVE_A070 16'hA070
`define TANH_LUT_NEGATIVE_A078 16'hA078
`define TANH_LUT_NEGATIVE_A080 16'hA080
`define TANH_LUT_NEGATIVE_A088 16'hA088
`define TANH_LUT_NEGATIVE_A090 16'hA090
`define TANH_LUT_NEGATIVE_A098 16'hA098
`define TANH_LUT_NEGATIVE_A0A0 16'hA0A0
`define TANH_LUT_NEGATIVE_A0A8 16'hA0A8
`define TANH_LUT_NEGATIVE_A0B0 16'hA0B0
`define TANH_LUT_NEGATIVE_A0B8 16'hA0B8
`define TANH_LUT_NEGATIVE_A0C0 16'hA0C0
`define TANH_LUT_NEGATIVE_A0C8 16'hA0C8
`define TANH_LUT_NEGATIVE_A0D0 16'hA0D0
`define TANH_LUT_NEGATIVE_A0D8 16'hA0D8
`define TANH_LUT_NEGATIVE_A0E0 16'hA0E0
`define TANH_LUT_NEGATIVE_A0E8 16'hA0E8
`define TANH_LUT_NEGATIVE_A0F0 16'hA0F0
`define TANH_LUT_NEGATIVE_A0F8 16'hA0F8
`define TANH_LUT_NEGATIVE_A100 16'hA100
`define TANH_LUT_NEGATIVE_A108 16'hA108
`define TANH_LUT_NEGATIVE_A110 16'hA110
`define TANH_LUT_NEGATIVE_A118 16'hA118
`define TANH_LUT_NEGATIVE_A120 16'hA120
`define TANH_LUT_NEGATIVE_A128 16'hA128
`define TANH_LUT_NEGATIVE_A130 16'hA130
`define TANH_LUT_NEGATIVE_A138 16'hA138
`define TANH_LUT_NEGATIVE_A140 16'hA140
`define TANH_LUT_NEGATIVE_A148 16'hA148
`define TANH_LUT_NEGATIVE_A150 16'hA150
`define TANH_LUT_NEGATIVE_A158 16'hA158
`define TANH_LUT_NEGATIVE_A160 16'hA160
`define TANH_LUT_NEGATIVE_A168 16'hA168
`define TANH_LUT_NEGATIVE_A170 16'hA170
`define TANH_LUT_NEGATIVE_A178 16'hA178
`define TANH_LUT_NEGATIVE_A180 16'hA180
`define TANH_LUT_NEGATIVE_A188 16'hA188
`define TANH_LUT_NEGATIVE_A190 16'hA190
`define TANH_LUT_NEGATIVE_A198 16'hA198
`define TANH_LUT_NEGATIVE_A1A0 16'hA1A0
`define TANH_LUT_NEGATIVE_A1A8 16'hA1A8
`define TANH_LUT_NEGATIVE_A1B0 16'hA1B0
`define TANH_LUT_NEGATIVE_A1B8 16'hA1B8
`define TANH_LUT_NEGATIVE_A1C0 16'hA1C0
`define TANH_LUT_NEGATIVE_A1C8 16'hA1C8
`define TANH_LUT_NEGATIVE_A1D0 16'hA1D0
`define TANH_LUT_NEGATIVE_A1D8 16'hA1D8
`define TANH_LUT_NEGATIVE_A1E0 16'hA1E0
`define TANH_LUT_NEGATIVE_A1E8 16'hA1E8
`define TANH_LUT_NEGATIVE_A1F0 16'hA1F0
`define TANH_LUT_NEGATIVE_A1F8 16'hA1F8
`define TANH_LUT_NEGATIVE_A200 16'hA200
`define TANH_LUT_NEGATIVE_A208 16'hA208
`define TANH_LUT_NEGATIVE_A210 16'hA210
`define TANH_LUT_NEGATIVE_A218 16'hA218
`define TANH_LUT_NEGATIVE_A220 16'hA220
`define TANH_LUT_NEGATIVE_A228 16'hA228
`define TANH_LUT_NEGATIVE_A230 16'hA230
`define TANH_LUT_NEGATIVE_A238 16'hA238
`define TANH_LUT_NEGATIVE_A240 16'hA240
`define TANH_LUT_NEGATIVE_A248 16'hA248
`define TANH_LUT_NEGATIVE_A250 16'hA250
`define TANH_LUT_NEGATIVE_A258 16'hA258
`define TANH_LUT_NEGATIVE_A260 16'hA260
`define TANH_LUT_NEGATIVE_A268 16'hA268
`define TANH_LUT_NEGATIVE_A270 16'hA270
`define TANH_LUT_NEGATIVE_A278 16'hA278
`define TANH_LUT_NEGATIVE_A280 16'hA280
`define TANH_LUT_NEGATIVE_A288 16'hA288
`define TANH_LUT_NEGATIVE_A290 16'hA290
`define TANH_LUT_NEGATIVE_A298 16'hA298
`define TANH_LUT_NEGATIVE_A2A0 16'hA2A0
`define TANH_LUT_NEGATIVE_A2A8 16'hA2A8
`define TANH_LUT_NEGATIVE_A2B0 16'hA2B0
`define TANH_LUT_NEGATIVE_A2B8 16'hA2B8
`define TANH_LUT_NEGATIVE_A2C0 16'hA2C0
`define TANH_LUT_NEGATIVE_A2C8 16'hA2C8
`define TANH_LUT_NEGATIVE_A2D0 16'hA2D0
`define TANH_LUT_NEGATIVE_A2D8 16'hA2D8
`define TANH_LUT_NEGATIVE_A2E0 16'hA2E0
`define TANH_LUT_NEGATIVE_A2E8 16'hA2E8
`define TANH_LUT_NEGATIVE_A2F0 16'hA2F0
`define TANH_LUT_NEGATIVE_A2F8 16'hA2F8
`define TANH_LUT_NEGATIVE_A300 16'hA300
`define TANH_LUT_NEGATIVE_A308 16'hA308
`define TANH_LUT_NEGATIVE_A310 16'hA310
`define TANH_LUT_NEGATIVE_A318 16'hA318
`define TANH_LUT_NEGATIVE_A320 16'hA320
`define TANH_LUT_NEGATIVE_A328 16'hA328
`define TANH_LUT_NEGATIVE_A330 16'hA330
`define TANH_LUT_NEGATIVE_A338 16'hA338
`define TANH_LUT_NEGATIVE_A340 16'hA340
`define TANH_LUT_NEGATIVE_A348 16'hA348
`define TANH_LUT_NEGATIVE_A350 16'hA350
`define TANH_LUT_NEGATIVE_A358 16'hA358
`define TANH_LUT_NEGATIVE_A360 16'hA360
`define TANH_LUT_NEGATIVE_A368 16'hA368
`define TANH_LUT_NEGATIVE_A370 16'hA370
`define TANH_LUT_NEGATIVE_A378 16'hA378
`define TANH_LUT_NEGATIVE_A380 16'hA380
`define TANH_LUT_NEGATIVE_A388 16'hA388
`define TANH_LUT_NEGATIVE_A390 16'hA390
`define TANH_LUT_NEGATIVE_A398 16'hA398
`define TANH_LUT_NEGATIVE_A3A0 16'hA3A0
`define TANH_LUT_NEGATIVE_A3A8 16'hA3A8
`define TANH_LUT_NEGATIVE_A3B0 16'hA3B0
`define TANH_LUT_NEGATIVE_A3B8 16'hA3B8
`define TANH_LUT_NEGATIVE_A3C0 16'hA3C0
`define TANH_LUT_NEGATIVE_A3C8 16'hA3C8
`define TANH_LUT_NEGATIVE_A3D0 16'hA3D0
`define TANH_LUT_NEGATIVE_A3D8 16'hA3D8
`define TANH_LUT_NEGATIVE_A3E0 16'hA3E0
`define TANH_LUT_NEGATIVE_A3E8 16'hA3E8
`define TANH_LUT_NEGATIVE_A3F0 16'hA3F0
`define TANH_LUT_NEGATIVE_A3F8 16'hA3F8
`define TANH_LUT_NEGATIVE_A400 16'hA400
`define TANH_LUT_NEGATIVE_A408 16'hA408
`define TANH_LUT_NEGATIVE_A410 16'hA410
`define TANH_LUT_NEGATIVE_A418 16'hA418
`define TANH_LUT_NEGATIVE_A420 16'hA420
`define TANH_LUT_NEGATIVE_A428 16'hA428
`define TANH_LUT_NEGATIVE_A430 16'hA430
`define TANH_LUT_NEGATIVE_A438 16'hA438
`define TANH_LUT_NEGATIVE_A440 16'hA440
`define TANH_LUT_NEGATIVE_A448 16'hA448
`define TANH_LUT_NEGATIVE_A450 16'hA450
`define TANH_LUT_NEGATIVE_A458 16'hA458
`define TANH_LUT_NEGATIVE_A460 16'hA460
`define TANH_LUT_NEGATIVE_A468 16'hA468
`define TANH_LUT_NEGATIVE_A470 16'hA470
`define TANH_LUT_NEGATIVE_A478 16'hA478
`define TANH_LUT_NEGATIVE_A480 16'hA480
`define TANH_LUT_NEGATIVE_A488 16'hA488
`define TANH_LUT_NEGATIVE_A490 16'hA490
`define TANH_LUT_NEGATIVE_A498 16'hA498
`define TANH_LUT_NEGATIVE_A4A0 16'hA4A0
`define TANH_LUT_NEGATIVE_A4A8 16'hA4A8
`define TANH_LUT_NEGATIVE_A4B0 16'hA4B0
`define TANH_LUT_NEGATIVE_A4B8 16'hA4B8
`define TANH_LUT_NEGATIVE_A4C0 16'hA4C0
`define TANH_LUT_NEGATIVE_A4C8 16'hA4C8
`define TANH_LUT_NEGATIVE_A4D0 16'hA4D0
`define TANH_LUT_NEGATIVE_A4D8 16'hA4D8
`define TANH_LUT_NEGATIVE_A4E0 16'hA4E0
`define TANH_LUT_NEGATIVE_A4E8 16'hA4E8
`define TANH_LUT_NEGATIVE_A4F0 16'hA4F0
`define TANH_LUT_NEGATIVE_A4F8 16'hA4F8
`define TANH_LUT_NEGATIVE_A500 16'hA500
`define TANH_LUT_NEGATIVE_A508 16'hA508
`define TANH_LUT_NEGATIVE_A510 16'hA510
`define TANH_LUT_NEGATIVE_A518 16'hA518
`define TANH_LUT_NEGATIVE_A520 16'hA520
`define TANH_LUT_NEGATIVE_A528 16'hA528
`define TANH_LUT_NEGATIVE_A530 16'hA530
`define TANH_LUT_NEGATIVE_A538 16'hA538
`define TANH_LUT_NEGATIVE_A540 16'hA540
`define TANH_LUT_NEGATIVE_A548 16'hA548
`define TANH_LUT_NEGATIVE_A550 16'hA550
`define TANH_LUT_NEGATIVE_A558 16'hA558
`define TANH_LUT_NEGATIVE_A560 16'hA560
`define TANH_LUT_NEGATIVE_A568 16'hA568
`define TANH_LUT_NEGATIVE_A570 16'hA570
`define TANH_LUT_NEGATIVE_A578 16'hA578
`define TANH_LUT_NEGATIVE_A580 16'hA580
`define TANH_LUT_NEGATIVE_A588 16'hA588
`define TANH_LUT_NEGATIVE_A590 16'hA590
`define TANH_LUT_NEGATIVE_A598 16'hA598
`define TANH_LUT_NEGATIVE_A5A0 16'hA5A0
`define TANH_LUT_NEGATIVE_A5A8 16'hA5A8
`define TANH_LUT_NEGATIVE_A5B0 16'hA5B0
`define TANH_LUT_NEGATIVE_A5B8 16'hA5B8
`define TANH_LUT_NEGATIVE_A5C0 16'hA5C0
`define TANH_LUT_NEGATIVE_A5C8 16'hA5C8
`define TANH_LUT_NEGATIVE_A5D0 16'hA5D0
`define TANH_LUT_NEGATIVE_A5D8 16'hA5D8
`define TANH_LUT_NEGATIVE_A5E0 16'hA5E0
`define TANH_LUT_NEGATIVE_A5E8 16'hA5E8
`define TANH_LUT_NEGATIVE_A5F0 16'hA5F0
`define TANH_LUT_NEGATIVE_A5F8 16'hA5F8
`define TANH_LUT_NEGATIVE_A600 16'hA600
`define TANH_LUT_NEGATIVE_A608 16'hA608
`define TANH_LUT_NEGATIVE_A610 16'hA610
`define TANH_LUT_NEGATIVE_A618 16'hA618
`define TANH_LUT_NEGATIVE_A620 16'hA620
`define TANH_LUT_NEGATIVE_A628 16'hA628
`define TANH_LUT_NEGATIVE_A630 16'hA630
`define TANH_LUT_NEGATIVE_A638 16'hA638
`define TANH_LUT_NEGATIVE_A640 16'hA640
`define TANH_LUT_NEGATIVE_A648 16'hA648
`define TANH_LUT_NEGATIVE_A650 16'hA650
`define TANH_LUT_NEGATIVE_A658 16'hA658
`define TANH_LUT_NEGATIVE_A660 16'hA660
`define TANH_LUT_NEGATIVE_A668 16'hA668
`define TANH_LUT_NEGATIVE_A670 16'hA670
`define TANH_LUT_NEGATIVE_A678 16'hA678
`define TANH_LUT_NEGATIVE_A680 16'hA680
`define TANH_LUT_NEGATIVE_A688 16'hA688
`define TANH_LUT_NEGATIVE_A690 16'hA690
`define TANH_LUT_NEGATIVE_A698 16'hA698
`define TANH_LUT_NEGATIVE_A6A0 16'hA6A0
`define TANH_LUT_NEGATIVE_A6A8 16'hA6A8
`define TANH_LUT_NEGATIVE_A6B0 16'hA6B0
`define TANH_LUT_NEGATIVE_A6B8 16'hA6B8
`define TANH_LUT_NEGATIVE_A6C0 16'hA6C0
`define TANH_LUT_NEGATIVE_A6C8 16'hA6C8
`define TANH_LUT_NEGATIVE_A6D0 16'hA6D0
`define TANH_LUT_NEGATIVE_A6D8 16'hA6D8
`define TANH_LUT_NEGATIVE_A6E0 16'hA6E0
`define TANH_LUT_NEGATIVE_A6E8 16'hA6E8
`define TANH_LUT_NEGATIVE_A6F0 16'hA6F0
`define TANH_LUT_NEGATIVE_A6F8 16'hA6F8
`define TANH_LUT_NEGATIVE_A700 16'hA700
`define TANH_LUT_NEGATIVE_A708 16'hA708
`define TANH_LUT_NEGATIVE_A710 16'hA710
`define TANH_LUT_NEGATIVE_A718 16'hA718
`define TANH_LUT_NEGATIVE_A720 16'hA720
`define TANH_LUT_NEGATIVE_A728 16'hA728
`define TANH_LUT_NEGATIVE_A730 16'hA730
`define TANH_LUT_NEGATIVE_A738 16'hA738
`define TANH_LUT_NEGATIVE_A740 16'hA740
`define TANH_LUT_NEGATIVE_A748 16'hA747
`define TANH_LUT_NEGATIVE_A750 16'hA74F
`define TANH_LUT_NEGATIVE_A758 16'hA757
`define TANH_LUT_NEGATIVE_A760 16'hA75F
`define TANH_LUT_NEGATIVE_A768 16'hA767
`define TANH_LUT_NEGATIVE_A770 16'hA76F
`define TANH_LUT_NEGATIVE_A778 16'hA777
`define TANH_LUT_NEGATIVE_A780 16'hA77F
`define TANH_LUT_NEGATIVE_A788 16'hA787
`define TANH_LUT_NEGATIVE_A790 16'hA78F
`define TANH_LUT_NEGATIVE_A798 16'hA797
`define TANH_LUT_NEGATIVE_A7A0 16'hA79F
`define TANH_LUT_NEGATIVE_A7A8 16'hA7A7
`define TANH_LUT_NEGATIVE_A7B0 16'hA7AF
`define TANH_LUT_NEGATIVE_A7B8 16'hA7B7
`define TANH_LUT_NEGATIVE_A7C0 16'hA7BF
`define TANH_LUT_NEGATIVE_A7C8 16'hA7C7
`define TANH_LUT_NEGATIVE_A7D0 16'hA7CF
`define TANH_LUT_NEGATIVE_A7D8 16'hA7D7
`define TANH_LUT_NEGATIVE_A7E0 16'hA7DF
`define TANH_LUT_NEGATIVE_A7E8 16'hA7E7
`define TANH_LUT_NEGATIVE_A7F0 16'hA7EF
`define TANH_LUT_NEGATIVE_A7F8 16'hA7F7
`define TANH_LUT_NEGATIVE_A800 16'hA7FF
`define TANH_LUT_NEGATIVE_A808 16'hA808
`define TANH_LUT_NEGATIVE_A810 16'hA810
`define TANH_LUT_NEGATIVE_A818 16'hA818
`define TANH_LUT_NEGATIVE_A820 16'hA820
`define TANH_LUT_NEGATIVE_A828 16'hA828
`define TANH_LUT_NEGATIVE_A830 16'hA830
`define TANH_LUT_NEGATIVE_A838 16'hA838
`define TANH_LUT_NEGATIVE_A840 16'hA840
`define TANH_LUT_NEGATIVE_A848 16'hA848
`define TANH_LUT_NEGATIVE_A850 16'hA850
`define TANH_LUT_NEGATIVE_A858 16'hA858
`define TANH_LUT_NEGATIVE_A860 16'hA860
`define TANH_LUT_NEGATIVE_A868 16'hA868
`define TANH_LUT_NEGATIVE_A870 16'hA870
`define TANH_LUT_NEGATIVE_A878 16'hA878
`define TANH_LUT_NEGATIVE_A880 16'hA880
`define TANH_LUT_NEGATIVE_A888 16'hA888
`define TANH_LUT_NEGATIVE_A890 16'hA890
`define TANH_LUT_NEGATIVE_A898 16'hA897
`define TANH_LUT_NEGATIVE_A8A0 16'hA89F
`define TANH_LUT_NEGATIVE_A8A8 16'hA8A7
`define TANH_LUT_NEGATIVE_A8B0 16'hA8AF
`define TANH_LUT_NEGATIVE_A8B8 16'hA8B7
`define TANH_LUT_NEGATIVE_A8C0 16'hA8BF
`define TANH_LUT_NEGATIVE_A8C8 16'hA8C7
`define TANH_LUT_NEGATIVE_A8D0 16'hA8CF
`define TANH_LUT_NEGATIVE_A8D8 16'hA8D7
`define TANH_LUT_NEGATIVE_A8E0 16'hA8DF
`define TANH_LUT_NEGATIVE_A8E8 16'hA8E7
`define TANH_LUT_NEGATIVE_A8F0 16'hA8EF
`define TANH_LUT_NEGATIVE_A8F8 16'hA8F7
`define TANH_LUT_NEGATIVE_A900 16'hA8FF
`define TANH_LUT_NEGATIVE_A908 16'hA907
`define TANH_LUT_NEGATIVE_A910 16'hA90F
`define TANH_LUT_NEGATIVE_A918 16'hA917
`define TANH_LUT_NEGATIVE_A920 16'hA91F
`define TANH_LUT_NEGATIVE_A928 16'hA927
`define TANH_LUT_NEGATIVE_A930 16'hA92F
`define TANH_LUT_NEGATIVE_A938 16'hA937
`define TANH_LUT_NEGATIVE_A940 16'hA93F
`define TANH_LUT_NEGATIVE_A948 16'hA947
`define TANH_LUT_NEGATIVE_A950 16'hA94F
`define TANH_LUT_NEGATIVE_A958 16'hA957
`define TANH_LUT_NEGATIVE_A960 16'hA95F
`define TANH_LUT_NEGATIVE_A968 16'hA967
`define TANH_LUT_NEGATIVE_A970 16'hA96F
`define TANH_LUT_NEGATIVE_A978 16'hA977
`define TANH_LUT_NEGATIVE_A980 16'hA97F
`define TANH_LUT_NEGATIVE_A988 16'hA987
`define TANH_LUT_NEGATIVE_A990 16'hA98F
`define TANH_LUT_NEGATIVE_A998 16'hA997
`define TANH_LUT_NEGATIVE_A9A0 16'hA99F
`define TANH_LUT_NEGATIVE_A9A8 16'hA9A7
`define TANH_LUT_NEGATIVE_A9B0 16'hA9AF
`define TANH_LUT_NEGATIVE_A9B8 16'hA9B7
`define TANH_LUT_NEGATIVE_A9C0 16'hA9BF
`define TANH_LUT_NEGATIVE_A9C8 16'hA9C7
`define TANH_LUT_NEGATIVE_A9D0 16'hA9CF
`define TANH_LUT_NEGATIVE_A9D8 16'hA9D7
`define TANH_LUT_NEGATIVE_A9E0 16'hA9DF
`define TANH_LUT_NEGATIVE_A9E8 16'hA9E7
`define TANH_LUT_NEGATIVE_A9F0 16'hA9EF
`define TANH_LUT_NEGATIVE_A9F8 16'hA9F7
`define TANH_LUT_NEGATIVE_AA00 16'hA9FF
`define TANH_LUT_NEGATIVE_AA08 16'hAA07
`define TANH_LUT_NEGATIVE_AA10 16'hAA0F
`define TANH_LUT_NEGATIVE_AA18 16'hAA17
`define TANH_LUT_NEGATIVE_AA20 16'hAA1F
`define TANH_LUT_NEGATIVE_AA28 16'hAA27
`define TANH_LUT_NEGATIVE_AA30 16'hAA2F
`define TANH_LUT_NEGATIVE_AA38 16'hAA37
`define TANH_LUT_NEGATIVE_AA40 16'hAA3F
`define TANH_LUT_NEGATIVE_AA48 16'hAA47
`define TANH_LUT_NEGATIVE_AA50 16'hAA4F
`define TANH_LUT_NEGATIVE_AA58 16'hAA57
`define TANH_LUT_NEGATIVE_AA60 16'hAA5F
`define TANH_LUT_NEGATIVE_AA68 16'hAA67
`define TANH_LUT_NEGATIVE_AA70 16'hAA6F
`define TANH_LUT_NEGATIVE_AA78 16'hAA77
`define TANH_LUT_NEGATIVE_AA80 16'hAA7F
`define TANH_LUT_NEGATIVE_AA88 16'hAA87
`define TANH_LUT_NEGATIVE_AA90 16'hAA8F
`define TANH_LUT_NEGATIVE_AA98 16'hAA97
`define TANH_LUT_NEGATIVE_AAA0 16'hAA9E
`define TANH_LUT_NEGATIVE_AAA8 16'hAAA6
`define TANH_LUT_NEGATIVE_AAB0 16'hAAAE
`define TANH_LUT_NEGATIVE_AAB8 16'hAAB6
`define TANH_LUT_NEGATIVE_AAC0 16'hAABE
`define TANH_LUT_NEGATIVE_AAC8 16'hAAC6
`define TANH_LUT_NEGATIVE_AAD0 16'hAACE
`define TANH_LUT_NEGATIVE_AAD8 16'hAAD6
`define TANH_LUT_NEGATIVE_AAE0 16'hAADE
`define TANH_LUT_NEGATIVE_AAE8 16'hAAE6
`define TANH_LUT_NEGATIVE_AAF0 16'hAAEE
`define TANH_LUT_NEGATIVE_AAF8 16'hAAF6
`define TANH_LUT_NEGATIVE_AB00 16'hAAFE
`define TANH_LUT_NEGATIVE_AB08 16'hAB06
`define TANH_LUT_NEGATIVE_AB10 16'hAB0E
`define TANH_LUT_NEGATIVE_AB18 16'hAB16
`define TANH_LUT_NEGATIVE_AB20 16'hAB1E
`define TANH_LUT_NEGATIVE_AB28 16'hAB26
`define TANH_LUT_NEGATIVE_AB30 16'hAB2E
`define TANH_LUT_NEGATIVE_AB38 16'hAB36
`define TANH_LUT_NEGATIVE_AB40 16'hAB3E
`define TANH_LUT_NEGATIVE_AB48 16'hAB46
`define TANH_LUT_NEGATIVE_AB50 16'hAB4E
`define TANH_LUT_NEGATIVE_AB58 16'hAB56
`define TANH_LUT_NEGATIVE_AB60 16'hAB5E
`define TANH_LUT_NEGATIVE_AB68 16'hAB66
`define TANH_LUT_NEGATIVE_AB70 16'hAB6E
`define TANH_LUT_NEGATIVE_AB78 16'hAB76
`define TANH_LUT_NEGATIVE_AB80 16'hAB7E
`define TANH_LUT_NEGATIVE_AB88 16'hAB86
`define TANH_LUT_NEGATIVE_AB90 16'hAB8E
`define TANH_LUT_NEGATIVE_AB98 16'hAB96
`define TANH_LUT_NEGATIVE_ABA0 16'hAB9E
`define TANH_LUT_NEGATIVE_ABA8 16'hABA6
`define TANH_LUT_NEGATIVE_ABB0 16'hABAE
`define TANH_LUT_NEGATIVE_ABB8 16'hABB6
`define TANH_LUT_NEGATIVE_ABC0 16'hABBE
`define TANH_LUT_NEGATIVE_ABC8 16'hABC6
`define TANH_LUT_NEGATIVE_ABD0 16'hABCE
`define TANH_LUT_NEGATIVE_ABD8 16'hABD5
`define TANH_LUT_NEGATIVE_ABE0 16'hABDD
`define TANH_LUT_NEGATIVE_ABE8 16'hABE5
`define TANH_LUT_NEGATIVE_ABF0 16'hABED
`define TANH_LUT_NEGATIVE_ABF8 16'hABF5
`define TANH_LUT_NEGATIVE_AC00 16'hABFD
`define TANH_LUT_NEGATIVE_AC08 16'hAC07
`define TANH_LUT_NEGATIVE_AC10 16'hAC0F
`define TANH_LUT_NEGATIVE_AC18 16'hAC17
`define TANH_LUT_NEGATIVE_AC20 16'hAC1F
`define TANH_LUT_NEGATIVE_AC28 16'hAC27
`define TANH_LUT_NEGATIVE_AC30 16'hAC2E
`define TANH_LUT_NEGATIVE_AC38 16'hAC36
`define TANH_LUT_NEGATIVE_AC40 16'hAC3E
`define TANH_LUT_NEGATIVE_AC48 16'hAC46
`define TANH_LUT_NEGATIVE_AC50 16'hAC4E
`define TANH_LUT_NEGATIVE_AC58 16'hAC56
`define TANH_LUT_NEGATIVE_AC60 16'hAC5E
`define TANH_LUT_NEGATIVE_AC68 16'hAC66
`define TANH_LUT_NEGATIVE_AC70 16'hAC6E
`define TANH_LUT_NEGATIVE_AC78 16'hAC76
`define TANH_LUT_NEGATIVE_AC80 16'hAC7E
`define TANH_LUT_NEGATIVE_AC88 16'hAC86
`define TANH_LUT_NEGATIVE_AC90 16'hAC8E
`define TANH_LUT_NEGATIVE_AC98 16'hAC96
`define TANH_LUT_NEGATIVE_ACA0 16'hAC9E
`define TANH_LUT_NEGATIVE_ACA8 16'hACA6
`define TANH_LUT_NEGATIVE_ACB0 16'hACAE
`define TANH_LUT_NEGATIVE_ACB8 16'hACB6
`define TANH_LUT_NEGATIVE_ACC0 16'hACBE
`define TANH_LUT_NEGATIVE_ACC8 16'hACC6
`define TANH_LUT_NEGATIVE_ACD0 16'hACCE
`define TANH_LUT_NEGATIVE_ACD8 16'hACD6
`define TANH_LUT_NEGATIVE_ACE0 16'hACDE
`define TANH_LUT_NEGATIVE_ACE8 16'hACE6
`define TANH_LUT_NEGATIVE_ACF0 16'hACED
`define TANH_LUT_NEGATIVE_ACF8 16'hACF5
`define TANH_LUT_NEGATIVE_AD00 16'hACFD
`define TANH_LUT_NEGATIVE_AD08 16'hAD05
`define TANH_LUT_NEGATIVE_AD10 16'hAD0D
`define TANH_LUT_NEGATIVE_AD18 16'hAD15
`define TANH_LUT_NEGATIVE_AD20 16'hAD1D
`define TANH_LUT_NEGATIVE_AD28 16'hAD25
`define TANH_LUT_NEGATIVE_AD30 16'hAD2D
`define TANH_LUT_NEGATIVE_AD38 16'hAD35
`define TANH_LUT_NEGATIVE_AD40 16'hAD3D
`define TANH_LUT_NEGATIVE_AD48 16'hAD45
`define TANH_LUT_NEGATIVE_AD50 16'hAD4D
`define TANH_LUT_NEGATIVE_AD58 16'hAD55
`define TANH_LUT_NEGATIVE_AD60 16'hAD5D
`define TANH_LUT_NEGATIVE_AD68 16'hAD65
`define TANH_LUT_NEGATIVE_AD70 16'hAD6D
`define TANH_LUT_NEGATIVE_AD78 16'hAD75
`define TANH_LUT_NEGATIVE_AD80 16'hAD7D
`define TANH_LUT_NEGATIVE_AD88 16'hAD84
`define TANH_LUT_NEGATIVE_AD90 16'hAD8C
`define TANH_LUT_NEGATIVE_AD98 16'hAD94
`define TANH_LUT_NEGATIVE_ADA0 16'hAD9C
`define TANH_LUT_NEGATIVE_ADA8 16'hADA4
`define TANH_LUT_NEGATIVE_ADB0 16'hADAC
`define TANH_LUT_NEGATIVE_ADB8 16'hADB4
`define TANH_LUT_NEGATIVE_ADC0 16'hADBC
`define TANH_LUT_NEGATIVE_ADC8 16'hADC4
`define TANH_LUT_NEGATIVE_ADD0 16'hADCC
`define TANH_LUT_NEGATIVE_ADD8 16'hADD4
`define TANH_LUT_NEGATIVE_ADE0 16'hADDC
`define TANH_LUT_NEGATIVE_ADE8 16'hADE4
`define TANH_LUT_NEGATIVE_ADF0 16'hADEC
`define TANH_LUT_NEGATIVE_ADF8 16'hADF4
`define TANH_LUT_NEGATIVE_AE00 16'hADFC
`define TANH_LUT_NEGATIVE_AE08 16'hAE03
`define TANH_LUT_NEGATIVE_AE10 16'hAE0B
`define TANH_LUT_NEGATIVE_AE18 16'hAE13
`define TANH_LUT_NEGATIVE_AE20 16'hAE1B
`define TANH_LUT_NEGATIVE_AE28 16'hAE23
`define TANH_LUT_NEGATIVE_AE30 16'hAE2B
`define TANH_LUT_NEGATIVE_AE38 16'hAE33
`define TANH_LUT_NEGATIVE_AE40 16'hAE3B
`define TANH_LUT_NEGATIVE_AE48 16'hAE43
`define TANH_LUT_NEGATIVE_AE50 16'hAE4B
`define TANH_LUT_NEGATIVE_AE58 16'hAE53
`define TANH_LUT_NEGATIVE_AE60 16'hAE5B
`define TANH_LUT_NEGATIVE_AE68 16'hAE63
`define TANH_LUT_NEGATIVE_AE70 16'hAE6A
`define TANH_LUT_NEGATIVE_AE78 16'hAE72
`define TANH_LUT_NEGATIVE_AE80 16'hAE7A
`define TANH_LUT_NEGATIVE_AE88 16'hAE82
`define TANH_LUT_NEGATIVE_AE90 16'hAE8A
`define TANH_LUT_NEGATIVE_AE98 16'hAE92
`define TANH_LUT_NEGATIVE_AEA0 16'hAE9A
`define TANH_LUT_NEGATIVE_AEA8 16'hAEA2
`define TANH_LUT_NEGATIVE_AEB0 16'hAEAA
`define TANH_LUT_NEGATIVE_AEB8 16'hAEB2
`define TANH_LUT_NEGATIVE_AEC0 16'hAEBA
`define TANH_LUT_NEGATIVE_AEC8 16'hAEC2
`define TANH_LUT_NEGATIVE_AED0 16'hAEC9
`define TANH_LUT_NEGATIVE_AED8 16'hAED1
`define TANH_LUT_NEGATIVE_AEE0 16'hAED9
`define TANH_LUT_NEGATIVE_AEE8 16'hAEE1
`define TANH_LUT_NEGATIVE_AEF0 16'hAEE9
`define TANH_LUT_NEGATIVE_AEF8 16'hAEF1
`define TANH_LUT_NEGATIVE_AF00 16'hAEF9
`define TANH_LUT_NEGATIVE_AF08 16'hAF01
`define TANH_LUT_NEGATIVE_AF10 16'hAF09
`define TANH_LUT_NEGATIVE_AF18 16'hAF11
`define TANH_LUT_NEGATIVE_AF20 16'hAF19
`define TANH_LUT_NEGATIVE_AF28 16'hAF20
`define TANH_LUT_NEGATIVE_AF30 16'hAF28
`define TANH_LUT_NEGATIVE_AF38 16'hAF30
`define TANH_LUT_NEGATIVE_AF40 16'hAF38
`define TANH_LUT_NEGATIVE_AF48 16'hAF40
`define TANH_LUT_NEGATIVE_AF50 16'hAF48
`define TANH_LUT_NEGATIVE_AF58 16'hAF50
`define TANH_LUT_NEGATIVE_AF60 16'hAF58
`define TANH_LUT_NEGATIVE_AF68 16'hAF60
`define TANH_LUT_NEGATIVE_AF70 16'hAF67
`define TANH_LUT_NEGATIVE_AF78 16'hAF6F
`define TANH_LUT_NEGATIVE_AF80 16'hAF77
`define TANH_LUT_NEGATIVE_AF88 16'hAF7F
`define TANH_LUT_NEGATIVE_AF90 16'hAF87
`define TANH_LUT_NEGATIVE_AF98 16'hAF8F
`define TANH_LUT_NEGATIVE_AFA0 16'hAF97
`define TANH_LUT_NEGATIVE_AFA8 16'hAF9F
`define TANH_LUT_NEGATIVE_AFB0 16'hAFA7
`define TANH_LUT_NEGATIVE_AFB8 16'hAFAE
`define TANH_LUT_NEGATIVE_AFC0 16'hAFB6
`define TANH_LUT_NEGATIVE_AFC8 16'hAFBE
`define TANH_LUT_NEGATIVE_AFD0 16'hAFC6
`define TANH_LUT_NEGATIVE_AFD8 16'hAFCE
`define TANH_LUT_NEGATIVE_AFE0 16'hAFD6
`define TANH_LUT_NEGATIVE_AFE8 16'hAFDE
`define TANH_LUT_NEGATIVE_AFF0 16'hAFE6
`define TANH_LUT_NEGATIVE_AFF8 16'hAFEE
`define TANH_LUT_NEGATIVE_B000 16'hAFF5
`define TANH_LUT_NEGATIVE_B008 16'hB003
`define TANH_LUT_NEGATIVE_B010 16'hB00A
`define TANH_LUT_NEGATIVE_B018 16'hB012
`define TANH_LUT_NEGATIVE_B020 16'hB01A
`define TANH_LUT_NEGATIVE_B028 16'hB022
`define TANH_LUT_NEGATIVE_B030 16'hB02A
`define TANH_LUT_NEGATIVE_B038 16'hB032
`define TANH_LUT_NEGATIVE_B040 16'hB03A
`define TANH_LUT_NEGATIVE_B048 16'hB042
`define TANH_LUT_NEGATIVE_B050 16'hB049
`define TANH_LUT_NEGATIVE_B058 16'hB051
`define TANH_LUT_NEGATIVE_B060 16'hB059
`define TANH_LUT_NEGATIVE_B068 16'hB061
`define TANH_LUT_NEGATIVE_B070 16'hB069
`define TANH_LUT_NEGATIVE_B078 16'hB071
`define TANH_LUT_NEGATIVE_B080 16'hB078
`define TANH_LUT_NEGATIVE_B088 16'hB080
`define TANH_LUT_NEGATIVE_B090 16'hB088
`define TANH_LUT_NEGATIVE_B098 16'hB090
`define TANH_LUT_NEGATIVE_B0A0 16'hB098
`define TANH_LUT_NEGATIVE_B0A8 16'hB0A0
`define TANH_LUT_NEGATIVE_B0B0 16'hB0A7
`define TANH_LUT_NEGATIVE_B0B8 16'hB0AF
`define TANH_LUT_NEGATIVE_B0C0 16'hB0B7
`define TANH_LUT_NEGATIVE_B0C8 16'hB0BF
`define TANH_LUT_NEGATIVE_B0D0 16'hB0C7
`define TANH_LUT_NEGATIVE_B0D8 16'hB0CF
`define TANH_LUT_NEGATIVE_B0E0 16'hB0D6
`define TANH_LUT_NEGATIVE_B0E8 16'hB0DE
`define TANH_LUT_NEGATIVE_B0F0 16'hB0E6
`define TANH_LUT_NEGATIVE_B0F8 16'hB0EE
`define TANH_LUT_NEGATIVE_B100 16'hB0F6
`define TANH_LUT_NEGATIVE_B108 16'hB0FD
`define TANH_LUT_NEGATIVE_B110 16'hB105
`define TANH_LUT_NEGATIVE_B118 16'hB10D
`define TANH_LUT_NEGATIVE_B120 16'hB115
`define TANH_LUT_NEGATIVE_B128 16'hB11D
`define TANH_LUT_NEGATIVE_B130 16'hB124
`define TANH_LUT_NEGATIVE_B138 16'hB12C
`define TANH_LUT_NEGATIVE_B140 16'hB134
`define TANH_LUT_NEGATIVE_B148 16'hB13C
`define TANH_LUT_NEGATIVE_B150 16'hB144
`define TANH_LUT_NEGATIVE_B158 16'hB14B
`define TANH_LUT_NEGATIVE_B160 16'hB153
`define TANH_LUT_NEGATIVE_B168 16'hB15B
`define TANH_LUT_NEGATIVE_B170 16'hB163
`define TANH_LUT_NEGATIVE_B178 16'hB16B
`define TANH_LUT_NEGATIVE_B180 16'hB172
`define TANH_LUT_NEGATIVE_B188 16'hB17A
`define TANH_LUT_NEGATIVE_B190 16'hB182
`define TANH_LUT_NEGATIVE_B198 16'hB18A
`define TANH_LUT_NEGATIVE_B1A0 16'hB191
`define TANH_LUT_NEGATIVE_B1A8 16'hB199
`define TANH_LUT_NEGATIVE_B1B0 16'hB1A1
`define TANH_LUT_NEGATIVE_B1B8 16'hB1A9
`define TANH_LUT_NEGATIVE_B1C0 16'hB1B0
`define TANH_LUT_NEGATIVE_B1C8 16'hB1B8
`define TANH_LUT_NEGATIVE_B1D0 16'hB1C0
`define TANH_LUT_NEGATIVE_B1D8 16'hB1C8
`define TANH_LUT_NEGATIVE_B1E0 16'hB1CF
`define TANH_LUT_NEGATIVE_B1E8 16'hB1D7
`define TANH_LUT_NEGATIVE_B1F0 16'hB1DF
`define TANH_LUT_NEGATIVE_B1F8 16'hB1E7
`define TANH_LUT_NEGATIVE_B200 16'hB1EE
`define TANH_LUT_NEGATIVE_B208 16'hB1F6
`define TANH_LUT_NEGATIVE_B210 16'hB1FE
`define TANH_LUT_NEGATIVE_B218 16'hB205
`define TANH_LUT_NEGATIVE_B220 16'hB20D
`define TANH_LUT_NEGATIVE_B228 16'hB215
`define TANH_LUT_NEGATIVE_B230 16'hB21D
`define TANH_LUT_NEGATIVE_B238 16'hB224
`define TANH_LUT_NEGATIVE_B240 16'hB22C
`define TANH_LUT_NEGATIVE_B248 16'hB234
`define TANH_LUT_NEGATIVE_B250 16'hB23B
`define TANH_LUT_NEGATIVE_B258 16'hB243
`define TANH_LUT_NEGATIVE_B260 16'hB24B
`define TANH_LUT_NEGATIVE_B268 16'hB252
`define TANH_LUT_NEGATIVE_B270 16'hB25A
`define TANH_LUT_NEGATIVE_B278 16'hB262
`define TANH_LUT_NEGATIVE_B280 16'hB269
`define TANH_LUT_NEGATIVE_B288 16'hB271
`define TANH_LUT_NEGATIVE_B290 16'hB279
`define TANH_LUT_NEGATIVE_B298 16'hB281
`define TANH_LUT_NEGATIVE_B2A0 16'hB288
`define TANH_LUT_NEGATIVE_B2A8 16'hB290
`define TANH_LUT_NEGATIVE_B2B0 16'hB298
`define TANH_LUT_NEGATIVE_B2B8 16'hB29F
`define TANH_LUT_NEGATIVE_B2C0 16'hB2A7
`define TANH_LUT_NEGATIVE_B2C8 16'hB2AE
`define TANH_LUT_NEGATIVE_B2D0 16'hB2B6
`define TANH_LUT_NEGATIVE_B2D8 16'hB2BE
`define TANH_LUT_NEGATIVE_B2E0 16'hB2C5
`define TANH_LUT_NEGATIVE_B2E8 16'hB2CD
`define TANH_LUT_NEGATIVE_B2F0 16'hB2D5
`define TANH_LUT_NEGATIVE_B2F8 16'hB2DC
`define TANH_LUT_NEGATIVE_B300 16'hB2E4
`define TANH_LUT_NEGATIVE_B308 16'hB2EC
`define TANH_LUT_NEGATIVE_B310 16'hB2F3
`define TANH_LUT_NEGATIVE_B318 16'hB2FB
`define TANH_LUT_NEGATIVE_B320 16'hB302
`define TANH_LUT_NEGATIVE_B328 16'hB30A
`define TANH_LUT_NEGATIVE_B330 16'hB312
`define TANH_LUT_NEGATIVE_B338 16'hB319
`define TANH_LUT_NEGATIVE_B340 16'hB321
`define TANH_LUT_NEGATIVE_B348 16'hB328
`define TANH_LUT_NEGATIVE_B350 16'hB330
`define TANH_LUT_NEGATIVE_B358 16'hB338
`define TANH_LUT_NEGATIVE_B360 16'hB33F
`define TANH_LUT_NEGATIVE_B368 16'hB347
`define TANH_LUT_NEGATIVE_B370 16'hB34E
`define TANH_LUT_NEGATIVE_B378 16'hB356
`define TANH_LUT_NEGATIVE_B380 16'hB35E
`define TANH_LUT_NEGATIVE_B388 16'hB365
`define TANH_LUT_NEGATIVE_B390 16'hB36D
`define TANH_LUT_NEGATIVE_B398 16'hB374
`define TANH_LUT_NEGATIVE_B3A0 16'hB37C
`define TANH_LUT_NEGATIVE_B3A8 16'hB383
`define TANH_LUT_NEGATIVE_B3B0 16'hB38B
`define TANH_LUT_NEGATIVE_B3B8 16'hB393
`define TANH_LUT_NEGATIVE_B3C0 16'hB39A
`define TANH_LUT_NEGATIVE_B3C8 16'hB3A2
`define TANH_LUT_NEGATIVE_B3D0 16'hB3A9
`define TANH_LUT_NEGATIVE_B3D8 16'hB3B1
`define TANH_LUT_NEGATIVE_B3E0 16'hB3B8
`define TANH_LUT_NEGATIVE_B3E8 16'hB3C0
`define TANH_LUT_NEGATIVE_B3F0 16'hB3C7
`define TANH_LUT_NEGATIVE_B3F8 16'hB3CF
`define TANH_LUT_NEGATIVE_B400 16'hB3D6
`define TANH_LUT_NEGATIVE_B408 16'hB3E5
`define TANH_LUT_NEGATIVE_B410 16'hB3F4
`define TANH_LUT_NEGATIVE_B418 16'hB402
`define TANH_LUT_NEGATIVE_B420 16'hB409
`define TANH_LUT_NEGATIVE_B428 16'hB411
`define TANH_LUT_NEGATIVE_B430 16'hB418
`define TANH_LUT_NEGATIVE_B438 16'hB420
`define TANH_LUT_NEGATIVE_B440 16'hB427
`define TANH_LUT_NEGATIVE_B448 16'hB42F
`define TANH_LUT_NEGATIVE_B450 16'hB436
`define TANH_LUT_NEGATIVE_B458 16'hB43D
`define TANH_LUT_NEGATIVE_B460 16'hB445
`define TANH_LUT_NEGATIVE_B468 16'hB44C
`define TANH_LUT_NEGATIVE_B470 16'hB454
`define TANH_LUT_NEGATIVE_B478 16'hB45B
`define TANH_LUT_NEGATIVE_B480 16'hB463
`define TANH_LUT_NEGATIVE_B488 16'hB46A
`define TANH_LUT_NEGATIVE_B490 16'hB471
`define TANH_LUT_NEGATIVE_B498 16'hB479
`define TANH_LUT_NEGATIVE_B4A0 16'hB480
`define TANH_LUT_NEGATIVE_B4A8 16'hB487
`define TANH_LUT_NEGATIVE_B4B0 16'hB48F
`define TANH_LUT_NEGATIVE_B4B8 16'hB496
`define TANH_LUT_NEGATIVE_B4C0 16'hB49D
`define TANH_LUT_NEGATIVE_B4C8 16'hB4A5
`define TANH_LUT_NEGATIVE_B4D0 16'hB4AC
`define TANH_LUT_NEGATIVE_B4D8 16'hB4B3
`define TANH_LUT_NEGATIVE_B4E0 16'hB4BB
`define TANH_LUT_NEGATIVE_B4E8 16'hB4C2
`define TANH_LUT_NEGATIVE_B4F0 16'hB4C9
`define TANH_LUT_NEGATIVE_B4F8 16'hB4D1
`define TANH_LUT_NEGATIVE_B500 16'hB4D8
`define TANH_LUT_NEGATIVE_B508 16'hB4DF
`define TANH_LUT_NEGATIVE_B510 16'hB4E6
`define TANH_LUT_NEGATIVE_B518 16'hB4EE
`define TANH_LUT_NEGATIVE_B520 16'hB4F5
`define TANH_LUT_NEGATIVE_B528 16'hB4FC
`define TANH_LUT_NEGATIVE_B530 16'hB503
`define TANH_LUT_NEGATIVE_B538 16'hB50B
`define TANH_LUT_NEGATIVE_B540 16'hB512
`define TANH_LUT_NEGATIVE_B548 16'hB519
`define TANH_LUT_NEGATIVE_B550 16'hB520
`define TANH_LUT_NEGATIVE_B558 16'hB527
`define TANH_LUT_NEGATIVE_B560 16'hB52E
`define TANH_LUT_NEGATIVE_B568 16'hB536
`define TANH_LUT_NEGATIVE_B570 16'hB53D
`define TANH_LUT_NEGATIVE_B578 16'hB544
`define TANH_LUT_NEGATIVE_B580 16'hB54B
`define TANH_LUT_NEGATIVE_B588 16'hB552
`define TANH_LUT_NEGATIVE_B590 16'hB559
`define TANH_LUT_NEGATIVE_B598 16'hB560
`define TANH_LUT_NEGATIVE_B5A0 16'hB567
`define TANH_LUT_NEGATIVE_B5A8 16'hB56F
`define TANH_LUT_NEGATIVE_B5B0 16'hB576
`define TANH_LUT_NEGATIVE_B5B8 16'hB57D
`define TANH_LUT_NEGATIVE_B5C0 16'hB584
`define TANH_LUT_NEGATIVE_B5C8 16'hB58B
`define TANH_LUT_NEGATIVE_B5D0 16'hB592
`define TANH_LUT_NEGATIVE_B5D8 16'hB599
`define TANH_LUT_NEGATIVE_B5E0 16'hB5A0
`define TANH_LUT_NEGATIVE_B5E8 16'hB5A7
`define TANH_LUT_NEGATIVE_B5F0 16'hB5AE
`define TANH_LUT_NEGATIVE_B5F8 16'hB5B5
`define TANH_LUT_NEGATIVE_B600 16'hB5BC
`define TANH_LUT_NEGATIVE_B608 16'hB5C3
`define TANH_LUT_NEGATIVE_B610 16'hB5CA
`define TANH_LUT_NEGATIVE_B618 16'hB5D1
`define TANH_LUT_NEGATIVE_B620 16'hB5D8
`define TANH_LUT_NEGATIVE_B628 16'hB5DF
`define TANH_LUT_NEGATIVE_B630 16'hB5E5
`define TANH_LUT_NEGATIVE_B638 16'hB5EC
`define TANH_LUT_NEGATIVE_B640 16'hB5F3
`define TANH_LUT_NEGATIVE_B648 16'hB5FA
`define TANH_LUT_NEGATIVE_B650 16'hB601
`define TANH_LUT_NEGATIVE_B658 16'hB608
`define TANH_LUT_NEGATIVE_B660 16'hB60F
`define TANH_LUT_NEGATIVE_B668 16'hB616
`define TANH_LUT_NEGATIVE_B670 16'hB61C
`define TANH_LUT_NEGATIVE_B678 16'hB623
`define TANH_LUT_NEGATIVE_B680 16'hB62A
`define TANH_LUT_NEGATIVE_B688 16'hB631
`define TANH_LUT_NEGATIVE_B690 16'hB638
`define TANH_LUT_NEGATIVE_B698 16'hB63F
`define TANH_LUT_NEGATIVE_B6A0 16'hB645
`define TANH_LUT_NEGATIVE_B6A8 16'hB64C
`define TANH_LUT_NEGATIVE_B6B0 16'hB653
`define TANH_LUT_NEGATIVE_B6B8 16'hB65A
`define TANH_LUT_NEGATIVE_B6C0 16'hB660
`define TANH_LUT_NEGATIVE_B6C8 16'hB667
`define TANH_LUT_NEGATIVE_B6D0 16'hB66E
`define TANH_LUT_NEGATIVE_B6D8 16'hB674
`define TANH_LUT_NEGATIVE_B6E0 16'hB67B
`define TANH_LUT_NEGATIVE_B6E8 16'hB682
`define TANH_LUT_NEGATIVE_B6F0 16'hB688
`define TANH_LUT_NEGATIVE_B6F8 16'hB68F
`define TANH_LUT_NEGATIVE_B700 16'hB696
`define TANH_LUT_NEGATIVE_B708 16'hB69C
`define TANH_LUT_NEGATIVE_B710 16'hB6A3
`define TANH_LUT_NEGATIVE_B718 16'hB6AA
`define TANH_LUT_NEGATIVE_B720 16'hB6B0
`define TANH_LUT_NEGATIVE_B728 16'hB6B7
`define TANH_LUT_NEGATIVE_B730 16'hB6BD
`define TANH_LUT_NEGATIVE_B738 16'hB6C4
`define TANH_LUT_NEGATIVE_B740 16'hB6CB
`define TANH_LUT_NEGATIVE_B748 16'hB6D1
`define TANH_LUT_NEGATIVE_B750 16'hB6D8
`define TANH_LUT_NEGATIVE_B758 16'hB6DE
`define TANH_LUT_NEGATIVE_B760 16'hB6E5
`define TANH_LUT_NEGATIVE_B768 16'hB6EB
`define TANH_LUT_NEGATIVE_B770 16'hB6F2
`define TANH_LUT_NEGATIVE_B778 16'hB6F8
`define TANH_LUT_NEGATIVE_B780 16'hB6FF
`define TANH_LUT_NEGATIVE_B788 16'hB705
`define TANH_LUT_NEGATIVE_B790 16'hB70C
`define TANH_LUT_NEGATIVE_B798 16'hB712
`define TANH_LUT_NEGATIVE_B7A0 16'hB719
`define TANH_LUT_NEGATIVE_B7A8 16'hB71F
`define TANH_LUT_NEGATIVE_B7B0 16'hB725
`define TANH_LUT_NEGATIVE_B7B8 16'hB72C
`define TANH_LUT_NEGATIVE_B7C0 16'hB732
`define TANH_LUT_NEGATIVE_B7C8 16'hB739
`define TANH_LUT_NEGATIVE_B7D0 16'hB73F
`define TANH_LUT_NEGATIVE_B7D8 16'hB745
`define TANH_LUT_NEGATIVE_B7E0 16'hB74C
`define TANH_LUT_NEGATIVE_B7E8 16'hB752
`define TANH_LUT_NEGATIVE_B7F0 16'hB758
`define TANH_LUT_NEGATIVE_B7F8 16'hB75F
`define TANH_LUT_NEGATIVE_B800 16'hB765
`define TANH_LUT_NEGATIVE_B808 16'hB771
`define TANH_LUT_NEGATIVE_B810 16'hB77E
`define TANH_LUT_NEGATIVE_B818 16'hB78A
`define TANH_LUT_NEGATIVE_B820 16'hB797
`define TANH_LUT_NEGATIVE_B828 16'hB7A3
`define TANH_LUT_NEGATIVE_B830 16'hB7B0
`define TANH_LUT_NEGATIVE_B838 16'hB7BC
`define TANH_LUT_NEGATIVE_B840 16'hB7C8
`define TANH_LUT_NEGATIVE_B848 16'hB7D4
`define TANH_LUT_NEGATIVE_B850 16'hB7E0
`define TANH_LUT_NEGATIVE_B858 16'hB7EC
`define TANH_LUT_NEGATIVE_B860 16'hB7F9
`define TANH_LUT_NEGATIVE_B868 16'hB802
`define TANH_LUT_NEGATIVE_B870 16'hB808
`define TANH_LUT_NEGATIVE_B878 16'hB80E
`define TANH_LUT_NEGATIVE_B880 16'hB814
`define TANH_LUT_NEGATIVE_B888 16'hB81A
`define TANH_LUT_NEGATIVE_B890 16'hB820
`define TANH_LUT_NEGATIVE_B898 16'hB826
`define TANH_LUT_NEGATIVE_B8A0 16'hB82C
`define TANH_LUT_NEGATIVE_B8A8 16'hB831
`define TANH_LUT_NEGATIVE_B8B0 16'hB837
`define TANH_LUT_NEGATIVE_B8B8 16'hB83D
`define TANH_LUT_NEGATIVE_B8C0 16'hB843
`define TANH_LUT_NEGATIVE_B8C8 16'hB848
`define TANH_LUT_NEGATIVE_B8D0 16'hB84E
`define TANH_LUT_NEGATIVE_B8D8 16'hB854
`define TANH_LUT_NEGATIVE_B8E0 16'hB859
`define TANH_LUT_NEGATIVE_B8E8 16'hB85F
`define TANH_LUT_NEGATIVE_B8F0 16'hB865
`define TANH_LUT_NEGATIVE_B8F8 16'hB86A
`define TANH_LUT_NEGATIVE_B900 16'hB870
`define TANH_LUT_NEGATIVE_B908 16'hB875
`define TANH_LUT_NEGATIVE_B910 16'hB87B
`define TANH_LUT_NEGATIVE_B918 16'hB880
`define TANH_LUT_NEGATIVE_B920 16'hB886
`define TANH_LUT_NEGATIVE_B928 16'hB88B
`define TANH_LUT_NEGATIVE_B930 16'hB891
`define TANH_LUT_NEGATIVE_B938 16'hB896
`define TANH_LUT_NEGATIVE_B940 16'hB89B
`define TANH_LUT_NEGATIVE_B948 16'hB8A1
`define TANH_LUT_NEGATIVE_B950 16'hB8A6
`define TANH_LUT_NEGATIVE_B958 16'hB8AB
`define TANH_LUT_NEGATIVE_B960 16'hB8B1
`define TANH_LUT_NEGATIVE_B968 16'hB8B6
`define TANH_LUT_NEGATIVE_B970 16'hB8BB
`define TANH_LUT_NEGATIVE_B978 16'hB8C0
`define TANH_LUT_NEGATIVE_B980 16'hB8C5
`define TANH_LUT_NEGATIVE_B988 16'hB8CB
`define TANH_LUT_NEGATIVE_B990 16'hB8D0
`define TANH_LUT_NEGATIVE_B998 16'hB8D5
`define TANH_LUT_NEGATIVE_B9A0 16'hB8DA
`define TANH_LUT_NEGATIVE_B9A8 16'hB8DF
`define TANH_LUT_NEGATIVE_B9B0 16'hB8E4
`define TANH_LUT_NEGATIVE_B9B8 16'hB8E9
`define TANH_LUT_NEGATIVE_B9C0 16'hB8EE
`define TANH_LUT_NEGATIVE_B9C8 16'hB8F3
`define TANH_LUT_NEGATIVE_B9D0 16'hB8F8
`define TANH_LUT_NEGATIVE_B9D8 16'hB8FD
`define TANH_LUT_NEGATIVE_B9E0 16'hB902
`define TANH_LUT_NEGATIVE_B9E8 16'hB906
`define TANH_LUT_NEGATIVE_B9F0 16'hB90B
`define TANH_LUT_NEGATIVE_B9F8 16'hB910
`define TANH_LUT_NEGATIVE_BA00 16'hB915
`define TANH_LUT_NEGATIVE_BA08 16'hB91A
`define TANH_LUT_NEGATIVE_BA10 16'hB91E
`define TANH_LUT_NEGATIVE_BA18 16'hB923
`define TANH_LUT_NEGATIVE_BA20 16'hB928
`define TANH_LUT_NEGATIVE_BA28 16'hB92C
`define TANH_LUT_NEGATIVE_BA30 16'hB931
`define TANH_LUT_NEGATIVE_BA38 16'hB936
`define TANH_LUT_NEGATIVE_BA40 16'hB93A
`define TANH_LUT_NEGATIVE_BA48 16'hB93F
`define TANH_LUT_NEGATIVE_BA50 16'hB943
`define TANH_LUT_NEGATIVE_BA58 16'hB948
`define TANH_LUT_NEGATIVE_BA60 16'hB94C
`define TANH_LUT_NEGATIVE_BA68 16'hB951
`define TANH_LUT_NEGATIVE_BA70 16'hB955
`define TANH_LUT_NEGATIVE_BA78 16'hB95A
`define TANH_LUT_NEGATIVE_BA80 16'hB95E
`define TANH_LUT_NEGATIVE_BA88 16'hB963
`define TANH_LUT_NEGATIVE_BA90 16'hB967
`define TANH_LUT_NEGATIVE_BA98 16'hB96B
`define TANH_LUT_NEGATIVE_BAA0 16'hB970
`define TANH_LUT_NEGATIVE_BAA8 16'hB974
`define TANH_LUT_NEGATIVE_BAB0 16'hB978
`define TANH_LUT_NEGATIVE_BAB8 16'hB97C
`define TANH_LUT_NEGATIVE_BAC0 16'hB981
`define TANH_LUT_NEGATIVE_BAC8 16'hB985
`define TANH_LUT_NEGATIVE_BAD0 16'hB989
`define TANH_LUT_NEGATIVE_BAD8 16'hB98D
`define TANH_LUT_NEGATIVE_BAE0 16'hB991
`define TANH_LUT_NEGATIVE_BAE8 16'hB995
`define TANH_LUT_NEGATIVE_BAF0 16'hB999
`define TANH_LUT_NEGATIVE_BAF8 16'hB99E
`define TANH_LUT_NEGATIVE_BB00 16'hB9A2
`define TANH_LUT_NEGATIVE_BB08 16'hB9A6
`define TANH_LUT_NEGATIVE_BB10 16'hB9AA
`define TANH_LUT_NEGATIVE_BB18 16'hB9AE
`define TANH_LUT_NEGATIVE_BB20 16'hB9B2
`define TANH_LUT_NEGATIVE_BB28 16'hB9B6
`define TANH_LUT_NEGATIVE_BB30 16'hB9B9
`define TANH_LUT_NEGATIVE_BB38 16'hB9BD
`define TANH_LUT_NEGATIVE_BB40 16'hB9C1
`define TANH_LUT_NEGATIVE_BB48 16'hB9C5
`define TANH_LUT_NEGATIVE_BB50 16'hB9C9
`define TANH_LUT_NEGATIVE_BB58 16'hB9CD
`define TANH_LUT_NEGATIVE_BB60 16'hB9D0
`define TANH_LUT_NEGATIVE_BB68 16'hB9D4
`define TANH_LUT_NEGATIVE_BB70 16'hB9D8
`define TANH_LUT_NEGATIVE_BB78 16'hB9DC
`define TANH_LUT_NEGATIVE_BB80 16'hB9DF
`define TANH_LUT_NEGATIVE_BB88 16'hB9E3
`define TANH_LUT_NEGATIVE_BB90 16'hB9E7
`define TANH_LUT_NEGATIVE_BB98 16'hB9EA
`define TANH_LUT_NEGATIVE_BBA0 16'hB9EE
`define TANH_LUT_NEGATIVE_BBA8 16'hB9F2
`define TANH_LUT_NEGATIVE_BBB0 16'hB9F5
`define TANH_LUT_NEGATIVE_BBB8 16'hB9F9
`define TANH_LUT_NEGATIVE_BBC0 16'hB9FC
`define TANH_LUT_NEGATIVE_BBC8 16'hBA00
`define TANH_LUT_NEGATIVE_BBD0 16'hBA03
`define TANH_LUT_NEGATIVE_BBD8 16'hBA07
`define TANH_LUT_NEGATIVE_BBE0 16'hBA0A
`define TANH_LUT_NEGATIVE_BBE8 16'hBA0E
`define TANH_LUT_NEGATIVE_BBF0 16'hBA11
`define TANH_LUT_NEGATIVE_BBF8 16'hBA14
`define TANH_LUT_NEGATIVE_BC00 16'hBA18
`define TANH_LUT_NEGATIVE_BC08 16'hBA1E
`define TANH_LUT_NEGATIVE_BC10 16'hBA25
`define TANH_LUT_NEGATIVE_BC18 16'hBA2C
`define TANH_LUT_NEGATIVE_BC20 16'hBA32
`define TANH_LUT_NEGATIVE_BC28 16'hBA38
`define TANH_LUT_NEGATIVE_BC30 16'hBA3F
`define TANH_LUT_NEGATIVE_BC38 16'hBA45
`define TANH_LUT_NEGATIVE_BC40 16'hBA4B
`define TANH_LUT_NEGATIVE_BC48 16'hBA51
`define TANH_LUT_NEGATIVE_BC50 16'hBA57
`define TANH_LUT_NEGATIVE_BC58 16'hBA5D
`define TANH_LUT_NEGATIVE_BC60 16'hBA63
`define TANH_LUT_NEGATIVE_BC68 16'hBA69
`define TANH_LUT_NEGATIVE_BC70 16'hBA6E
`define TANH_LUT_NEGATIVE_BC78 16'hBA74
`define TANH_LUT_NEGATIVE_BC80 16'hBA79
`define TANH_LUT_NEGATIVE_BC88 16'hBA7F
`define TANH_LUT_NEGATIVE_BC90 16'hBA84
`define TANH_LUT_NEGATIVE_BC98 16'hBA8A
`define TANH_LUT_NEGATIVE_BCA0 16'hBA8F
`define TANH_LUT_NEGATIVE_BCA8 16'hBA94
`define TANH_LUT_NEGATIVE_BCB0 16'hBA99
`define TANH_LUT_NEGATIVE_BCB8 16'hBA9E
`define TANH_LUT_NEGATIVE_BCC0 16'hBAA3
`define TANH_LUT_NEGATIVE_BCC8 16'hBAA8
`define TANH_LUT_NEGATIVE_BCD0 16'hBAAD
`define TANH_LUT_NEGATIVE_BCD8 16'hBAB2
`define TANH_LUT_NEGATIVE_BCE0 16'hBAB7
`define TANH_LUT_NEGATIVE_BCE8 16'hBABC
`define TANH_LUT_NEGATIVE_BCF0 16'hBAC0
`define TANH_LUT_NEGATIVE_BCF8 16'hBAC5
`define TANH_LUT_NEGATIVE_BD00 16'hBAC9
`define TANH_LUT_NEGATIVE_BD08 16'hBACE
`define TANH_LUT_NEGATIVE_BD10 16'hBAD2
`define TANH_LUT_NEGATIVE_BD18 16'hBAD6
`define TANH_LUT_NEGATIVE_BD20 16'hBADB
`define TANH_LUT_NEGATIVE_BD28 16'hBADF
`define TANH_LUT_NEGATIVE_BD30 16'hBAE3
`define TANH_LUT_NEGATIVE_BD38 16'hBAE7
`define TANH_LUT_NEGATIVE_BD40 16'hBAEB
`define TANH_LUT_NEGATIVE_BD48 16'hBAEF
`define TANH_LUT_NEGATIVE_BD50 16'hBAF3
`define TANH_LUT_NEGATIVE_BD58 16'hBAF7
`define TANH_LUT_NEGATIVE_BD60 16'hBAFB
`define TANH_LUT_NEGATIVE_BD68 16'hBAFF
`define TANH_LUT_NEGATIVE_BD70 16'hBB03
`define TANH_LUT_NEGATIVE_BD78 16'hBB06
`define TANH_LUT_NEGATIVE_BD80 16'hBB0A
`define TANH_LUT_NEGATIVE_BD88 16'hBB0D
`define TANH_LUT_NEGATIVE_BD90 16'hBB11
`define TANH_LUT_NEGATIVE_BD98 16'hBB15
`define TANH_LUT_NEGATIVE_BDA0 16'hBB18
`define TANH_LUT_NEGATIVE_BDA8 16'hBB1B
`define TANH_LUT_NEGATIVE_BDB0 16'hBB1F
`define TANH_LUT_NEGATIVE_BDB8 16'hBB22
`define TANH_LUT_NEGATIVE_BDC0 16'hBB25
`define TANH_LUT_NEGATIVE_BDC8 16'hBB28
`define TANH_LUT_NEGATIVE_BDD0 16'hBB2C
`define TANH_LUT_NEGATIVE_BDD8 16'hBB2F
`define TANH_LUT_NEGATIVE_BDE0 16'hBB32
`define TANH_LUT_NEGATIVE_BDE8 16'hBB35
`define TANH_LUT_NEGATIVE_BDF0 16'hBB38
`define TANH_LUT_NEGATIVE_BDF8 16'hBB3B
`define TANH_LUT_NEGATIVE_BE00 16'hBB3E
`define TANH_LUT_NEGATIVE_BE08 16'hBB41
`define TANH_LUT_NEGATIVE_BE10 16'hBB43
`define TANH_LUT_NEGATIVE_BE18 16'hBB46
`define TANH_LUT_NEGATIVE_BE20 16'hBB49
`define TANH_LUT_NEGATIVE_BE28 16'hBB4C
`define TANH_LUT_NEGATIVE_BE30 16'hBB4E
`define TANH_LUT_NEGATIVE_BE38 16'hBB51
`define TANH_LUT_NEGATIVE_BE40 16'hBB54
`define TANH_LUT_NEGATIVE_BE48 16'hBB56
`define TANH_LUT_NEGATIVE_BE50 16'hBB59
`define TANH_LUT_NEGATIVE_BE58 16'hBB5B
`define TANH_LUT_NEGATIVE_BE60 16'hBB5E
`define TANH_LUT_NEGATIVE_BE68 16'hBB60
`define TANH_LUT_NEGATIVE_BE70 16'hBB62
`define TANH_LUT_NEGATIVE_BE78 16'hBB65
`define TANH_LUT_NEGATIVE_BE80 16'hBB67
`define TANH_LUT_NEGATIVE_BE88 16'hBB69
`define TANH_LUT_NEGATIVE_BE90 16'hBB6C
`define TANH_LUT_NEGATIVE_BE98 16'hBB6E
`define TANH_LUT_NEGATIVE_BEA0 16'hBB70
`define TANH_LUT_NEGATIVE_BEA8 16'hBB72
`define TANH_LUT_NEGATIVE_BEB0 16'hBB74
`define TANH_LUT_NEGATIVE_BEB8 16'hBB76
`define TANH_LUT_NEGATIVE_BEC0 16'hBB78
`define TANH_LUT_NEGATIVE_BEC8 16'hBB7B
`define TANH_LUT_NEGATIVE_BED0 16'hBB7D
`define TANH_LUT_NEGATIVE_BED8 16'hBB7E
`define TANH_LUT_NEGATIVE_BEE0 16'hBB80
`define TANH_LUT_NEGATIVE_BEE8 16'hBB82
`define TANH_LUT_NEGATIVE_BEF0 16'hBB84
`define TANH_LUT_NEGATIVE_BEF8 16'hBB86
`define TANH_LUT_NEGATIVE_BF00 16'hBB88
`define TANH_LUT_NEGATIVE_BF08 16'hBB8A
`define TANH_LUT_NEGATIVE_BF10 16'hBB8C
`define TANH_LUT_NEGATIVE_BF18 16'hBB8D
`define TANH_LUT_NEGATIVE_BF20 16'hBB8F
`define TANH_LUT_NEGATIVE_BF28 16'hBB91
`define TANH_LUT_NEGATIVE_BF30 16'hBB92
`define TANH_LUT_NEGATIVE_BF38 16'hBB94
`define TANH_LUT_NEGATIVE_BF40 16'hBB96
`define TANH_LUT_NEGATIVE_BF48 16'hBB97
`define TANH_LUT_NEGATIVE_BF50 16'hBB99
`define TANH_LUT_NEGATIVE_BF58 16'hBB9A
`define TANH_LUT_NEGATIVE_BF60 16'hBB9C
`define TANH_LUT_NEGATIVE_BF68 16'hBB9D
`define TANH_LUT_NEGATIVE_BF70 16'hBB9F
`define TANH_LUT_NEGATIVE_BF78 16'hBBA0
`define TANH_LUT_NEGATIVE_BF80 16'hBBA2
`define TANH_LUT_NEGATIVE_BF88 16'hBBA3
`define TANH_LUT_NEGATIVE_BF90 16'hBBA5
`define TANH_LUT_NEGATIVE_BF98 16'hBBA6
`define TANH_LUT_NEGATIVE_BFA0 16'hBBA7
`define TANH_LUT_NEGATIVE_BFA8 16'hBBA9
`define TANH_LUT_NEGATIVE_BFB0 16'hBBAA
`define TANH_LUT_NEGATIVE_BFB8 16'hBBAB
`define TANH_LUT_NEGATIVE_BFC0 16'hBBAD
`define TANH_LUT_NEGATIVE_BFC8 16'hBBAE
`define TANH_LUT_NEGATIVE_BFD0 16'hBBAF
`define TANH_LUT_NEGATIVE_BFD8 16'hBBB0
`define TANH_LUT_NEGATIVE_BFE0 16'hBBB2
`define TANH_LUT_NEGATIVE_BFE8 16'hBBB3
`define TANH_LUT_NEGATIVE_BFF0 16'hBBB4
`define TANH_LUT_NEGATIVE_BFF8 16'hBBB5
`define TANH_LUT_NEGATIVE_C000 16'hBBB6
`define TANH_LUT_NEGATIVE_C008 16'hBBB9
`define TANH_LUT_NEGATIVE_C010 16'hBBBB
`define TANH_LUT_NEGATIVE_C018 16'hBBBD
`define TANH_LUT_NEGATIVE_C020 16'hBBBF
`define TANH_LUT_NEGATIVE_C028 16'hBBC1
`define TANH_LUT_NEGATIVE_C030 16'hBBC3
`define TANH_LUT_NEGATIVE_C038 16'hBBC5
`define TANH_LUT_NEGATIVE_C040 16'hBBC6
`define TANH_LUT_NEGATIVE_C048 16'hBBC8
`define TANH_LUT_NEGATIVE_C050 16'hBBCA
`define TANH_LUT_NEGATIVE_C058 16'hBBCB
`define TANH_LUT_NEGATIVE_C060 16'hBBCD
`define TANH_LUT_NEGATIVE_C068 16'hBBCF
`define TANH_LUT_NEGATIVE_C070 16'hBBD0
`define TANH_LUT_NEGATIVE_C078 16'hBBD2
`define TANH_LUT_NEGATIVE_C080 16'hBBD3
`define TANH_LUT_NEGATIVE_C088 16'hBBD4
`define TANH_LUT_NEGATIVE_C090 16'hBBD6
`define TANH_LUT_NEGATIVE_C098 16'hBBD7
`define TANH_LUT_NEGATIVE_C0A0 16'hBBD8
`define TANH_LUT_NEGATIVE_C0A8 16'hBBD9
`define TANH_LUT_NEGATIVE_C0B0 16'hBBDB
`define TANH_LUT_NEGATIVE_C0B8 16'hBBDC
`define TANH_LUT_NEGATIVE_C0C0 16'hBBDD
`define TANH_LUT_NEGATIVE_C0C8 16'hBBDE
`define TANH_LUT_NEGATIVE_C0D0 16'hBBDF
`define TANH_LUT_NEGATIVE_C0D8 16'hBBE0
`define TANH_LUT_NEGATIVE_C0E0 16'hBBE1
`define TANH_LUT_NEGATIVE_C0E8 16'hBBE2
`define TANH_LUT_NEGATIVE_C0F0 16'hBBE3
`define TANH_LUT_NEGATIVE_C0F8 16'hBBE4
`define TANH_LUT_NEGATIVE_C100 16'hBBE5
`define TANH_LUT_NEGATIVE_C108 16'hBBE5
`define TANH_LUT_NEGATIVE_C110 16'hBBE6
`define TANH_LUT_NEGATIVE_C118 16'hBBE7
`define TANH_LUT_NEGATIVE_C120 16'hBBE8
`define TANH_LUT_NEGATIVE_C128 16'hBBE9
`define TANH_LUT_NEGATIVE_C130 16'hBBE9
`define TANH_LUT_NEGATIVE_C138 16'hBBEA
`define TANH_LUT_NEGATIVE_C140 16'hBBEB
`define TANH_LUT_NEGATIVE_C148 16'hBBEB
`define TANH_LUT_NEGATIVE_C150 16'hBBEC
`define TANH_LUT_NEGATIVE_C158 16'hBBED
`define TANH_LUT_NEGATIVE_C160 16'hBBED
`define TANH_LUT_NEGATIVE_C168 16'hBBEE
`define TANH_LUT_NEGATIVE_C170 16'hBBEE
`define TANH_LUT_NEGATIVE_C178 16'hBBEF
`define TANH_LUT_NEGATIVE_C180 16'hBBEF
`define TANH_LUT_NEGATIVE_C188 16'hBBF0
`define TANH_LUT_NEGATIVE_C190 16'hBBF0
`define TANH_LUT_NEGATIVE_C198 16'hBBF1
`define TANH_LUT_NEGATIVE_C1A0 16'hBBF1
`define TANH_LUT_NEGATIVE_C1A8 16'hBBF2
`define TANH_LUT_NEGATIVE_C1B0 16'hBBF2
`define TANH_LUT_NEGATIVE_C1B8 16'hBBF3
`define TANH_LUT_NEGATIVE_C1C0 16'hBBF3
`define TANH_LUT_NEGATIVE_C1C8 16'hBBF3
`define TANH_LUT_NEGATIVE_C1D0 16'hBBF4
`define TANH_LUT_NEGATIVE_C1D8 16'hBBF4
`define TANH_LUT_NEGATIVE_C1E0 16'hBBF5
`define TANH_LUT_NEGATIVE_C1E8 16'hBBF5
`define TANH_LUT_NEGATIVE_C1F0 16'hBBF5
`define TANH_LUT_NEGATIVE_C1F8 16'hBBF6
`define TANH_LUT_NEGATIVE_C200 16'hBBF6
`define TANH_LUT_NEGATIVE_C208 16'hBBF6
`define TANH_LUT_NEGATIVE_C210 16'hBBF6
`define TANH_LUT_NEGATIVE_C218 16'hBBF7
`define TANH_LUT_NEGATIVE_C220 16'hBBF7
`define TANH_LUT_NEGATIVE_C228 16'hBBF7
`define TANH_LUT_NEGATIVE_C230 16'hBBF8
`define TANH_LUT_NEGATIVE_C238 16'hBBF8
`define TANH_LUT_NEGATIVE_C240 16'hBBF8
`define TANH_LUT_NEGATIVE_C248 16'hBBF8
`define TANH_LUT_NEGATIVE_C250 16'hBBF9
`define TANH_LUT_NEGATIVE_C258 16'hBBF9
`define TANH_LUT_NEGATIVE_C260 16'hBBF9
`define TANH_LUT_NEGATIVE_C268 16'hBBF9
`define TANH_LUT_NEGATIVE_C270 16'hBBF9
`define TANH_LUT_NEGATIVE_C278 16'hBBFA
`define TANH_LUT_NEGATIVE_C280 16'hBBFA
`define TANH_LUT_NEGATIVE_C288 16'hBBFA
`define TANH_LUT_NEGATIVE_C290 16'hBBFA
`define TANH_LUT_NEGATIVE_C298 16'hBBFA
`define TANH_LUT_NEGATIVE_C2A0 16'hBBFB
`define TANH_LUT_NEGATIVE_C2A8 16'hBBFB
`define TANH_LUT_NEGATIVE_C2B0 16'hBBFB
`define TANH_LUT_NEGATIVE_C2B8 16'hBBFB
`define TANH_LUT_NEGATIVE_C2C0 16'hBBFB
`define TANH_LUT_NEGATIVE_C2C8 16'hBBFB
`define TANH_LUT_NEGATIVE_C2D0 16'hBBFB
`define TANH_LUT_NEGATIVE_C2D8 16'hBBFC
