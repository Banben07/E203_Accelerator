`define CUBE_LUT_SIZE 1024
`define CUBE_LUT_BITS 10
`define CUBE_LUT_0 16'h1101010000000000
`define CUBE_LUT_1 16'h1101001111110100
`define CUBE_LUT_2 16'h1101001111101000
`define CUBE_LUT_3 16'h1101001111011100
`define CUBE_LUT_4 16'h1101001111010000
`define CUBE_LUT_5 16'h1101001111000101
`define CUBE_LUT_6 16'h1101001110111001
`define CUBE_LUT_7 16'h1101001110101101
`define CUBE_LUT_8 16'h1101001110100001
`define CUBE_LUT_9 16'h1101001110010110
`define CUBE_LUT_10 16'h1101001110001010
`define CUBE_LUT_11 16'h1101001101111111
`define CUBE_LUT_12 16'h1101001101110011
`define CUBE_LUT_13 16'h1101001101101000
`define CUBE_LUT_14 16'h1101001101011100
`define CUBE_LUT_15 16'h1101001101010001
`define CUBE_LUT_16 16'h1101001101000110
`define CUBE_LUT_17 16'h1101001100111011
`define CUBE_LUT_18 16'h1101001100101111
`define CUBE_LUT_19 16'h1101001100100100
`define CUBE_LUT_20 16'h1101001100011001
`define CUBE_LUT_21 16'h1101001100001110
`define CUBE_LUT_22 16'h1101001100000011
`define CUBE_LUT_23 16'h1101001011111000
`define CUBE_LUT_24 16'h1101001011101101
`define CUBE_LUT_25 16'h1101001011100010
`define CUBE_LUT_26 16'h1101001011010111
`define CUBE_LUT_27 16'h1101001011001101
`define CUBE_LUT_28 16'h1101001011000010
`define CUBE_LUT_29 16'h1101001010110111
`define CUBE_LUT_30 16'h1101001010101100
`define CUBE_LUT_31 16'h1101001010100010
`define CUBE_LUT_32 16'h1101001010010111
`define CUBE_LUT_33 16'h1101001010001101
`define CUBE_LUT_34 16'h1101001010000010
`define CUBE_LUT_35 16'h1101001001111000
`define CUBE_LUT_36 16'h1101001001101101
`define CUBE_LUT_37 16'h1101001001100011
`define CUBE_LUT_38 16'h1101001001011001
`define CUBE_LUT_39 16'h1101001001001110
`define CUBE_LUT_40 16'h1101001001000100
`define CUBE_LUT_41 16'h1101001000111010
`define CUBE_LUT_42 16'h1101001000110000
`define CUBE_LUT_43 16'h1101001000100110
`define CUBE_LUT_44 16'h1101001000011100
`define CUBE_LUT_45 16'h1101001000010010
`define CUBE_LUT_46 16'h1101001000001000
`define CUBE_LUT_47 16'h1101000111111110
`define CUBE_LUT_48 16'h1101000111110100
`define CUBE_LUT_49 16'h1101000111101010
`define CUBE_LUT_50 16'h1101000111100000
`define CUBE_LUT_51 16'h1101000111010110
`define CUBE_LUT_52 16'h1101000111001101
`define CUBE_LUT_53 16'h1101000111000011
`define CUBE_LUT_54 16'h1101000110111001
`define CUBE_LUT_55 16'h1101000110110000
`define CUBE_LUT_56 16'h1101000110100110
`define CUBE_LUT_57 16'h1101000110011101
`define CUBE_LUT_58 16'h1101000110010011
`define CUBE_LUT_59 16'h1101000110001010
`define CUBE_LUT_60 16'h1101000110000001
`define CUBE_LUT_61 16'h1101000101110111
`define CUBE_LUT_62 16'h1101000101101110
`define CUBE_LUT_63 16'h1101000101100101
`define CUBE_LUT_64 16'h1101000101011011
`define CUBE_LUT_65 16'h1101000101010010
`define CUBE_LUT_66 16'h1101000101001001
`define CUBE_LUT_67 16'h1101000101000000
`define CUBE_LUT_68 16'h1101000100110111
`define CUBE_LUT_69 16'h1101000100101110
`define CUBE_LUT_70 16'h1101000100100101
`define CUBE_LUT_71 16'h1101000100011100
`define CUBE_LUT_72 16'h1101000100010011
`define CUBE_LUT_73 16'h1101000100001010
`define CUBE_LUT_74 16'h1101000100000010
`define CUBE_LUT_75 16'h1101000011111001
`define CUBE_LUT_76 16'h1101000011110000
`define CUBE_LUT_77 16'h1101000011100111
`define CUBE_LUT_78 16'h1101000011011111
`define CUBE_LUT_79 16'h1101000011010110
`define CUBE_LUT_80 16'h1101000011001110
`define CUBE_LUT_81 16'h1101000011000101
`define CUBE_LUT_82 16'h1101000010111101
`define CUBE_LUT_83 16'h1101000010110100
`define CUBE_LUT_84 16'h1101000010101100
`define CUBE_LUT_85 16'h1101000010100011
`define CUBE_LUT_86 16'h1101000010011011
`define CUBE_LUT_87 16'h1101000010010011
`define CUBE_LUT_88 16'h1101000010001010
`define CUBE_LUT_89 16'h1101000010000010
`define CUBE_LUT_90 16'h1101000001111010
`define CUBE_LUT_91 16'h1101000001110010
`define CUBE_LUT_92 16'h1101000001101010
`define CUBE_LUT_93 16'h1101000001100010
`define CUBE_LUT_94 16'h1101000001011010
`define CUBE_LUT_95 16'h1101000001010010
`define CUBE_LUT_96 16'h1101000001001010
`define CUBE_LUT_97 16'h1101000001000010
`define CUBE_LUT_98 16'h1101000000111010
`define CUBE_LUT_99 16'h1101000000110010
`define CUBE_LUT_100 16'h1101000000101010
`define CUBE_LUT_101 16'h1101000000100011
`define CUBE_LUT_102 16'h1101000000011011
`define CUBE_LUT_103 16'h1101000000010011
`define CUBE_LUT_104 16'h1101000000001100
`define CUBE_LUT_105 16'h1101000000000100
`define CUBE_LUT_106 16'h1100111111111001
`define CUBE_LUT_107 16'h1100111111101010
`define CUBE_LUT_108 16'h1100111111011011
`define CUBE_LUT_109 16'h1100111111001100
`define CUBE_LUT_110 16'h1100111110111101
`define CUBE_LUT_111 16'h1100111110101110
`define CUBE_LUT_112 16'h1100111110100000
`define CUBE_LUT_113 16'h1100111110010001
`define CUBE_LUT_114 16'h1100111110000010
`define CUBE_LUT_115 16'h1100111101110100
`define CUBE_LUT_116 16'h1100111101100101
`define CUBE_LUT_117 16'h1100111101010111
`define CUBE_LUT_118 16'h1100111101001001
`define CUBE_LUT_119 16'h1100111100111011
`define CUBE_LUT_120 16'h1100111100101101
`define CUBE_LUT_121 16'h1100111100011111
`define CUBE_LUT_122 16'h1100111100010001
`define CUBE_LUT_123 16'h1100111100000011
`define CUBE_LUT_124 16'h1100111011110101
`define CUBE_LUT_125 16'h1100111011100111
`define CUBE_LUT_126 16'h1100111011011001
`define CUBE_LUT_127 16'h1100111011001100
`define CUBE_LUT_128 16'h1100111010111110
`define CUBE_LUT_129 16'h1100111010110001
`define CUBE_LUT_130 16'h1100111010100011
`define CUBE_LUT_131 16'h1100111010010110
`define CUBE_LUT_132 16'h1100111010001001
`define CUBE_LUT_133 16'h1100111001111100
`define CUBE_LUT_134 16'h1100111001101111
`define CUBE_LUT_135 16'h1100111001100001
`define CUBE_LUT_136 16'h1100111001010101
`define CUBE_LUT_137 16'h1100111001001000
`define CUBE_LUT_138 16'h1100111000111011
`define CUBE_LUT_139 16'h1100111000101110
`define CUBE_LUT_140 16'h1100111000100001
`define CUBE_LUT_141 16'h1100111000010101
`define CUBE_LUT_142 16'h1100111000001000
`define CUBE_LUT_143 16'h1100110111111100
`define CUBE_LUT_144 16'h1100110111101111
`define CUBE_LUT_145 16'h1100110111100011
`define CUBE_LUT_146 16'h1100110111010110
`define CUBE_LUT_147 16'h1100110111001010
`define CUBE_LUT_148 16'h1100110110111110
`define CUBE_LUT_149 16'h1100110110110010
`define CUBE_LUT_150 16'h1100110110100110
`define CUBE_LUT_151 16'h1100110110011010
`define CUBE_LUT_152 16'h1100110110001110
`define CUBE_LUT_153 16'h1100110110000010
`define CUBE_LUT_154 16'h1100110101110110
`define CUBE_LUT_155 16'h1100110101101011
`define CUBE_LUT_156 16'h1100110101011111
`define CUBE_LUT_157 16'h1100110101010100
`define CUBE_LUT_158 16'h1100110101001000
`define CUBE_LUT_159 16'h1100110100111101
`define CUBE_LUT_160 16'h1100110100110001
`define CUBE_LUT_161 16'h1100110100100110
`define CUBE_LUT_162 16'h1100110100011011
`define CUBE_LUT_163 16'h1100110100001111
`define CUBE_LUT_164 16'h1100110100000100
`define CUBE_LUT_165 16'h1100110011111001
`define CUBE_LUT_166 16'h1100110011101110
`define CUBE_LUT_167 16'h1100110011100011
`define CUBE_LUT_168 16'h1100110011011001
`define CUBE_LUT_169 16'h1100110011001110
`define CUBE_LUT_170 16'h1100110011000011
`define CUBE_LUT_171 16'h1100110010111000
`define CUBE_LUT_172 16'h1100110010101110
`define CUBE_LUT_173 16'h1100110010100011
`define CUBE_LUT_174 16'h1100110010011001
`define CUBE_LUT_175 16'h1100110010001110
`define CUBE_LUT_176 16'h1100110010000100
`define CUBE_LUT_177 16'h1100110001111010
`define CUBE_LUT_178 16'h1100110001101111
`define CUBE_LUT_179 16'h1100110001100101
`define CUBE_LUT_180 16'h1100110001011011
`define CUBE_LUT_181 16'h1100110001010001
`define CUBE_LUT_182 16'h1100110001000111
`define CUBE_LUT_183 16'h1100110000111101
`define CUBE_LUT_184 16'h1100110000110011
`define CUBE_LUT_185 16'h1100110000101001
`define CUBE_LUT_186 16'h1100110000100000
`define CUBE_LUT_187 16'h1100110000010110
`define CUBE_LUT_188 16'h1100110000001100
`define CUBE_LUT_189 16'h1100110000000011
`define CUBE_LUT_190 16'h1100101111110010
`define CUBE_LUT_191 16'h1100101111011111
`define CUBE_LUT_192 16'h1100101111001100
`define CUBE_LUT_193 16'h1100101110111010
`define CUBE_LUT_194 16'h1100101110100111
`define CUBE_LUT_195 16'h1100101110010101
`define CUBE_LUT_196 16'h1100101110000010
`define CUBE_LUT_197 16'h1100101101110000
`define CUBE_LUT_198 16'h1100101101011110
`define CUBE_LUT_199 16'h1100101101001100
`define CUBE_LUT_200 16'h1100101100111010
`define CUBE_LUT_201 16'h1100101100101000
`define CUBE_LUT_202 16'h1100101100010111
`define CUBE_LUT_203 16'h1100101100000101
`define CUBE_LUT_204 16'h1100101011110100
`define CUBE_LUT_205 16'h1100101011100011
`define CUBE_LUT_206 16'h1100101011010001
`define CUBE_LUT_207 16'h1100101011000000
`define CUBE_LUT_208 16'h1100101010101111
`define CUBE_LUT_209 16'h1100101010011110
`define CUBE_LUT_210 16'h1100101010001110
`define CUBE_LUT_211 16'h1100101001111101
`define CUBE_LUT_212 16'h1100101001101101
`define CUBE_LUT_213 16'h1100101001011100
`define CUBE_LUT_214 16'h1100101001001100
`define CUBE_LUT_215 16'h1100101000111100
`define CUBE_LUT_216 16'h1100101000101100
`define CUBE_LUT_217 16'h1100101000011100
`define CUBE_LUT_218 16'h1100101000001100
`define CUBE_LUT_219 16'h1100100111111100
`define CUBE_LUT_220 16'h1100100111101100
`define CUBE_LUT_221 16'h1100100111011101
`define CUBE_LUT_222 16'h1100100111001101
`define CUBE_LUT_223 16'h1100100110111110
`define CUBE_LUT_224 16'h1100100110101111
`define CUBE_LUT_225 16'h1100100110100000
`define CUBE_LUT_226 16'h1100100110010001
`define CUBE_LUT_227 16'h1100100110000010
`define CUBE_LUT_228 16'h1100100101110011
`define CUBE_LUT_229 16'h1100100101100100
`define CUBE_LUT_230 16'h1100100101010101
`define CUBE_LUT_231 16'h1100100101000111
`define CUBE_LUT_232 16'h1100100100111001
`define CUBE_LUT_233 16'h1100100100101010
`define CUBE_LUT_234 16'h1100100100011100
`define CUBE_LUT_235 16'h1100100100001110
`define CUBE_LUT_236 16'h1100100100000000
`define CUBE_LUT_237 16'h1100100011110010
`define CUBE_LUT_238 16'h1100100011100100
`define CUBE_LUT_239 16'h1100100011010111
`define CUBE_LUT_240 16'h1100100011001001
`define CUBE_LUT_241 16'h1100100010111100
`define CUBE_LUT_242 16'h1100100010101110
`define CUBE_LUT_243 16'h1100100010100001
`define CUBE_LUT_244 16'h1100100010010100
`define CUBE_LUT_245 16'h1100100010000111
`define CUBE_LUT_246 16'h1100100001111010
`define CUBE_LUT_247 16'h1100100001101101
`define CUBE_LUT_248 16'h1100100001100000
`define CUBE_LUT_249 16'h1100100001010011
`define CUBE_LUT_250 16'h1100100001000111
`define CUBE_LUT_251 16'h1100100000111010
`define CUBE_LUT_252 16'h1100100000101110
`define CUBE_LUT_253 16'h1100100000100001
`define CUBE_LUT_254 16'h1100100000010101
`define CUBE_LUT_255 16'h1100100000001001
`define CUBE_LUT_256 16'h1100011111111010
`define CUBE_LUT_257 16'h1100011111100010
`define CUBE_LUT_258 16'h1100011111001010
`define CUBE_LUT_259 16'h1100011110110011
`define CUBE_LUT_260 16'h1100011110011100
`define CUBE_LUT_261 16'h1100011110000100
`define CUBE_LUT_262 16'h1100011101101101
`define CUBE_LUT_263 16'h1100011101010111
`define CUBE_LUT_264 16'h1100011101000000
`define CUBE_LUT_265 16'h1100011100101010
`define CUBE_LUT_266 16'h1100011100010011
`define CUBE_LUT_267 16'h1100011011111101
`define CUBE_LUT_268 16'h1100011011101000
`define CUBE_LUT_269 16'h1100011011010010
`define CUBE_LUT_270 16'h1100011010111100
`define CUBE_LUT_271 16'h1100011010100111
`define CUBE_LUT_272 16'h1100011010010010
`define CUBE_LUT_273 16'h1100011001111101
`define CUBE_LUT_274 16'h1100011001101000
`define CUBE_LUT_275 16'h1100011001010011
`define CUBE_LUT_276 16'h1100011000111111
`define CUBE_LUT_277 16'h1100011000101011
`define CUBE_LUT_278 16'h1100011000010111
`define CUBE_LUT_279 16'h1100011000000011
`define CUBE_LUT_280 16'h1100010111101111
`define CUBE_LUT_281 16'h1100010111011011
`define CUBE_LUT_282 16'h1100010111001000
`define CUBE_LUT_283 16'h1100010110110101
`define CUBE_LUT_284 16'h1100010110100010
`define CUBE_LUT_285 16'h1100010110001111
`define CUBE_LUT_286 16'h1100010101111100
`define CUBE_LUT_287 16'h1100010101101001
`define CUBE_LUT_288 16'h1100010101010111
`define CUBE_LUT_289 16'h1100010101000101
`define CUBE_LUT_290 16'h1100010100110010
`define CUBE_LUT_291 16'h1100010100100001
`define CUBE_LUT_292 16'h1100010100001111
`define CUBE_LUT_293 16'h1100010011111101
`define CUBE_LUT_294 16'h1100010011101100
`define CUBE_LUT_295 16'h1100010011011010
`define CUBE_LUT_296 16'h1100010011001001
`define CUBE_LUT_297 16'h1100010010111000
`define CUBE_LUT_298 16'h1100010010100111
`define CUBE_LUT_299 16'h1100010010010111
`define CUBE_LUT_300 16'h1100010010000110
`define CUBE_LUT_301 16'h1100010001110110
`define CUBE_LUT_302 16'h1100010001100110
`define CUBE_LUT_303 16'h1100010001010110
`define CUBE_LUT_304 16'h1100010001000110
`define CUBE_LUT_305 16'h1100010000110110
`define CUBE_LUT_306 16'h1100010000100110
`define CUBE_LUT_307 16'h1100010000010111
`define CUBE_LUT_308 16'h1100010000001000
`define CUBE_LUT_309 16'h1100001111110001
`define CUBE_LUT_310 16'h1100001111010011
`define CUBE_LUT_311 16'h1100001110110110
`define CUBE_LUT_312 16'h1100001110011000
`define CUBE_LUT_313 16'h1100001101111011
`define CUBE_LUT_314 16'h1100001101011110
`define CUBE_LUT_315 16'h1100001101000010
`define CUBE_LUT_316 16'h1100001100100110
`define CUBE_LUT_317 16'h1100001100001010
`define CUBE_LUT_318 16'h1100001011101110
`define CUBE_LUT_319 16'h1100001011010011
`define CUBE_LUT_320 16'h1100001010111000
`define CUBE_LUT_321 16'h1100001010011101
`define CUBE_LUT_322 16'h1100001010000010
`define CUBE_LUT_323 16'h1100001001101000
`define CUBE_LUT_324 16'h1100001001001110
`define CUBE_LUT_325 16'h1100001000110100
`define CUBE_LUT_326 16'h1100001000011011
`define CUBE_LUT_327 16'h1100001000000010
`define CUBE_LUT_328 16'h1100000111101001
`define CUBE_LUT_329 16'h1100000111010000
`define CUBE_LUT_330 16'h1100000110111000
`define CUBE_LUT_331 16'h1100000110100000
`define CUBE_LUT_332 16'h1100000110001000
`define CUBE_LUT_333 16'h1100000101110001
`define CUBE_LUT_334 16'h1100000101011001
`define CUBE_LUT_335 16'h1100000101000010
`define CUBE_LUT_336 16'h1100000100101100
`define CUBE_LUT_337 16'h1100000100010101
`define CUBE_LUT_338 16'h1100000011111111
`define CUBE_LUT_339 16'h1100000011101001
`define CUBE_LUT_340 16'h1100000011010011
`define CUBE_LUT_341 16'h1100000010111110
`define CUBE_LUT_342 16'h1100000010101000
`define CUBE_LUT_343 16'h1100000010010011
`define CUBE_LUT_344 16'h1100000001111111
`define CUBE_LUT_345 16'h1100000001101010
`define CUBE_LUT_346 16'h1100000001010110
`define CUBE_LUT_347 16'h1100000001000010
`define CUBE_LUT_348 16'h1100000000101110
`define CUBE_LUT_349 16'h1100000000011011
`define CUBE_LUT_350 16'h1100000000000111
`define CUBE_LUT_351 16'h1011111111101001
`define CUBE_LUT_352 16'h1011111111000011
`define CUBE_LUT_353 16'h1011111110011110
`define CUBE_LUT_354 16'h1011111101111001
`define CUBE_LUT_355 16'h1011111101010101
`define CUBE_LUT_356 16'h1011111100110001
`define CUBE_LUT_357 16'h1011111100001110
`define CUBE_LUT_358 16'h1011111011101011
`define CUBE_LUT_359 16'h1011111011001001
`define CUBE_LUT_360 16'h1011111010100111
`define CUBE_LUT_361 16'h1011111010000101
`define CUBE_LUT_362 16'h1011111001100100
`define CUBE_LUT_363 16'h1011111001000100
`define CUBE_LUT_364 16'h1011111000100100
`define CUBE_LUT_365 16'h1011111000000100
`define CUBE_LUT_366 16'h1011110111100100
`define CUBE_LUT_367 16'h1011110111000110
`define CUBE_LUT_368 16'h1011110110100111
`define CUBE_LUT_369 16'h1011110110001001
`define CUBE_LUT_370 16'h1011110101101011
`define CUBE_LUT_371 16'h1011110101001110
`define CUBE_LUT_372 16'h1011110100110001
`define CUBE_LUT_373 16'h1011110100010101
`define CUBE_LUT_374 16'h1011110011111001
`define CUBE_LUT_375 16'h1011110011011101
`define CUBE_LUT_376 16'h1011110011000010
`define CUBE_LUT_377 16'h1011110010101000
`define CUBE_LUT_378 16'h1011110010001101
`define CUBE_LUT_379 16'h1011110001110011
`define CUBE_LUT_380 16'h1011110001011010
`define CUBE_LUT_381 16'h1011110001000000
`define CUBE_LUT_382 16'h1011110000101000
`define CUBE_LUT_383 16'h1011110000001111
`define CUBE_LUT_384 16'h1011101111101110
`define CUBE_LUT_385 16'h1011101110111111
`define CUBE_LUT_386 16'h1011101110010000
`define CUBE_LUT_387 16'h1011101101100010
`define CUBE_LUT_388 16'h1011101100110101
`define CUBE_LUT_389 16'h1011101100001000
`define CUBE_LUT_390 16'h1011101011011101
`define CUBE_LUT_391 16'h1011101010110010
`define CUBE_LUT_392 16'h1011101010000111
`define CUBE_LUT_393 16'h1011101001011110
`define CUBE_LUT_394 16'h1011101000110101
`define CUBE_LUT_395 16'h1011101000001101
`define CUBE_LUT_396 16'h1011100111100101
`define CUBE_LUT_397 16'h1011100110111110
`define CUBE_LUT_398 16'h1011100110011000
`define CUBE_LUT_399 16'h1011100101110011
`define CUBE_LUT_400 16'h1011100101001110
`define CUBE_LUT_401 16'h1011100100101001
`define CUBE_LUT_402 16'h1011100100000110
`define CUBE_LUT_403 16'h1011100011100011
`define CUBE_LUT_404 16'h1011100011000001
`define CUBE_LUT_405 16'h1011100010011111
`define CUBE_LUT_406 16'h1011100001111110
`define CUBE_LUT_407 16'h1011100001011110
`define CUBE_LUT_408 16'h1011100000111110
`define CUBE_LUT_409 16'h1011100000011111
`define CUBE_LUT_410 16'h1011100000000000
`define CUBE_LUT_411 16'h1011011111000100
`define CUBE_LUT_412 16'h1011011110001010
`define CUBE_LUT_413 16'h1011011101010000
`define CUBE_LUT_414 16'h1011011100011000
`define CUBE_LUT_415 16'h1011011011100000
`define CUBE_LUT_416 16'h1011011010101010
`define CUBE_LUT_417 16'h1011011001110101
`define CUBE_LUT_418 16'h1011011001000001
`define CUBE_LUT_419 16'h1011011000001110
`define CUBE_LUT_420 16'h1011010111011101
`define CUBE_LUT_421 16'h1011010110101100
`define CUBE_LUT_422 16'h1011010101111100
`define CUBE_LUT_423 16'h1011010101001110
`define CUBE_LUT_424 16'h1011010100100000
`define CUBE_LUT_425 16'h1011010011110100
`define CUBE_LUT_426 16'h1011010011001000
`define CUBE_LUT_427 16'h1011010010011110
`define CUBE_LUT_428 16'h1011010001110100
`define CUBE_LUT_429 16'h1011010001001100
`define CUBE_LUT_430 16'h1011010000100100
`define CUBE_LUT_431 16'h1011001111111100
`define CUBE_LUT_432 16'h1011001110110000
`define CUBE_LUT_433 16'h1011001101100111
`define CUBE_LUT_434 16'h1011001100100000
`define CUBE_LUT_435 16'h1011001011011010
`define CUBE_LUT_436 16'h1011001010010110
`define CUBE_LUT_437 16'h1011001001010100
`define CUBE_LUT_438 16'h1011001000010100
`define CUBE_LUT_439 16'h1011000111010101
`define CUBE_LUT_440 16'h1011000110011000
`define CUBE_LUT_441 16'h1011000101011101
`define CUBE_LUT_442 16'h1011000100100011
`define CUBE_LUT_443 16'h1011000011101011
`define CUBE_LUT_444 16'h1011000010110101
`define CUBE_LUT_445 16'h1011000010000000
`define CUBE_LUT_446 16'h1011000001001101
`define CUBE_LUT_447 16'h1011000000011011
`define CUBE_LUT_448 16'h1010111111010110
`define CUBE_LUT_449 16'h1010111101111001
`define CUBE_LUT_450 16'h1010111100011111
`define CUBE_LUT_451 16'h1010111011000111
`define CUBE_LUT_452 16'h1010111001110010
`define CUBE_LUT_453 16'h1010111000100001
`define CUBE_LUT_454 16'h1010110111010010
`define CUBE_LUT_455 16'h1010110110000101
`define CUBE_LUT_456 16'h1010110100111011
`define CUBE_LUT_457 16'h1010110011110100
`define CUBE_LUT_458 16'h1010110010110000
`define CUBE_LUT_459 16'h1010110001101110
`define CUBE_LUT_460 16'h1010110000101110
`define CUBE_LUT_461 16'h1010101111100010
`define CUBE_LUT_462 16'h1010101101101101
`define CUBE_LUT_463 16'h1010101011111100
`define CUBE_LUT_464 16'h1010101010001111
`define CUBE_LUT_465 16'h1010101000101000
`define CUBE_LUT_466 16'h1010100111000100
`define CUBE_LUT_467 16'h1010100101100101
`define CUBE_LUT_468 16'h1010100100001010
`define CUBE_LUT_469 16'h1010100010110011
`define CUBE_LUT_470 16'h1010100001100000
`define CUBE_LUT_471 16'h1010100000010001
`define CUBE_LUT_472 16'h1010011110001100
`define CUBE_LUT_473 16'h1010011011111101
`define CUBE_LUT_474 16'h1010011001110101
`define CUBE_LUT_475 16'h1010010111110100
`define CUBE_LUT_476 16'h1010010101111010
`define CUBE_LUT_477 16'h1010010100000111
`define CUBE_LUT_478 16'h1010010010011010
`define CUBE_LUT_479 16'h1010010000110100
`define CUBE_LUT_480 16'h1010001110100111
`define CUBE_LUT_481 16'h1010001011110010
`define CUBE_LUT_482 16'h1010001001001001
`define CUBE_LUT_483 16'h1010000110101011
`define CUBE_LUT_484 16'h1010000100011000
`define CUBE_LUT_485 16'h1010000010001111
`define CUBE_LUT_486 16'h1010000000001111
`define CUBE_LUT_487 16'h1001111100110100
`define CUBE_LUT_488 16'h1001111001011011
`define CUBE_LUT_489 16'h1001110110010100
`define CUBE_LUT_490 16'h1001110011011110
`define CUBE_LUT_491 16'h1001110000111000
`define CUBE_LUT_492 16'h1001101101000011
`define CUBE_LUT_493 16'h1001101000110100
`define CUBE_LUT_494 16'h1001100101000000
`define CUBE_LUT_495 16'h1001100001100110
`define CUBE_LUT_496 16'h1001011101001011
`define CUBE_LUT_497 16'h1001010111111001
`define CUBE_LUT_498 16'h1001010011010010
`define CUBE_LUT_499 16'h1001001110100111
`define CUBE_LUT_500 16'h1001000111110101
`define CUBE_LUT_501 16'h1001000010001001
`define CUBE_LUT_502 16'h1000111010111000
`define CUBE_LUT_503 16'h1000110011010000
`define CUBE_LUT_504 16'h1000101010011100
`define CUBE_LUT_505 16'h1000100001001110
`define CUBE_LUT_506 16'h1000010100110111
`define CUBE_LUT_507 16'h1000001011011011
`define CUBE_LUT_508 16'h1000000101011000
`define CUBE_LUT_509 16'h1000000001111101
`define CUBE_LUT_510 16'h1000000000011011
`define CUBE_LUT_511 16'h1000000000000001
`define CUBE_LUT_512 16'h0000000000000001
`define CUBE_LUT_513 16'h0000000000011011
`define CUBE_LUT_514 16'h0000000001111101
`define CUBE_LUT_515 16'h0000000101011000
`define CUBE_LUT_516 16'h0000001011011011
`define CUBE_LUT_517 16'h0000010100110111
`define CUBE_LUT_518 16'h0000100001001110
`define CUBE_LUT_519 16'h0000101010011100
`define CUBE_LUT_520 16'h0000110011010000
`define CUBE_LUT_521 16'h0000111010111000
`define CUBE_LUT_522 16'h0001000010001001
`define CUBE_LUT_523 16'h0001000111110101
`define CUBE_LUT_524 16'h0001001110100111
`define CUBE_LUT_525 16'h0001010011010010
`define CUBE_LUT_526 16'h0001010111111001
`define CUBE_LUT_527 16'h0001011101001011
`define CUBE_LUT_528 16'h0001100001100110
`define CUBE_LUT_529 16'h0001100101000000
`define CUBE_LUT_530 16'h0001101000110100
`define CUBE_LUT_531 16'h0001101101000011
`define CUBE_LUT_532 16'h0001110000111000
`define CUBE_LUT_533 16'h0001110011011110
`define CUBE_LUT_534 16'h0001110110010100
`define CUBE_LUT_535 16'h0001111001011011
`define CUBE_LUT_536 16'h0001111100110100
`define CUBE_LUT_537 16'h0010000000001111
`define CUBE_LUT_538 16'h0010000010001111
`define CUBE_LUT_539 16'h0010000100011000
`define CUBE_LUT_540 16'h0010000110101011
`define CUBE_LUT_541 16'h0010001001001001
`define CUBE_LUT_542 16'h0010001011110010
`define CUBE_LUT_543 16'h0010001110100111
`define CUBE_LUT_544 16'h0010010000110100
`define CUBE_LUT_545 16'h0010010010011010
`define CUBE_LUT_546 16'h0010010100000111
`define CUBE_LUT_547 16'h0010010101111010
`define CUBE_LUT_548 16'h0010010111110100
`define CUBE_LUT_549 16'h0010011001110101
`define CUBE_LUT_550 16'h0010011011111101
`define CUBE_LUT_551 16'h0010011110001100
`define CUBE_LUT_552 16'h0010100000010001
`define CUBE_LUT_553 16'h0010100001100000
`define CUBE_LUT_554 16'h0010100010110011
`define CUBE_LUT_555 16'h0010100100001010
`define CUBE_LUT_556 16'h0010100101100101
`define CUBE_LUT_557 16'h0010100111000100
`define CUBE_LUT_558 16'h0010101000101000
`define CUBE_LUT_559 16'h0010101010001111
`define CUBE_LUT_560 16'h0010101011111100
`define CUBE_LUT_561 16'h0010101101101101
`define CUBE_LUT_562 16'h0010101111100010
`define CUBE_LUT_563 16'h0010110000101110
`define CUBE_LUT_564 16'h0010110001101110
`define CUBE_LUT_565 16'h0010110010110000
`define CUBE_LUT_566 16'h0010110011110100
`define CUBE_LUT_567 16'h0010110100111011
`define CUBE_LUT_568 16'h0010110110000101
`define CUBE_LUT_569 16'h0010110111010010
`define CUBE_LUT_570 16'h0010111000100001
`define CUBE_LUT_571 16'h0010111001110010
`define CUBE_LUT_572 16'h0010111011000111
`define CUBE_LUT_573 16'h0010111100011111
`define CUBE_LUT_574 16'h0010111101111001
`define CUBE_LUT_575 16'h0010111111010110
`define CUBE_LUT_576 16'h0011000000011011
`define CUBE_LUT_577 16'h0011000001001101
`define CUBE_LUT_578 16'h0011000010000000
`define CUBE_LUT_579 16'h0011000010110101
`define CUBE_LUT_580 16'h0011000011101011
`define CUBE_LUT_581 16'h0011000100100011
`define CUBE_LUT_582 16'h0011000101011101
`define CUBE_LUT_583 16'h0011000110011000
`define CUBE_LUT_584 16'h0011000111010101
`define CUBE_LUT_585 16'h0011001000010100
`define CUBE_LUT_586 16'h0011001001010100
`define CUBE_LUT_587 16'h0011001010010110
`define CUBE_LUT_588 16'h0011001011011010
`define CUBE_LUT_589 16'h0011001100100000
`define CUBE_LUT_590 16'h0011001101100111
`define CUBE_LUT_591 16'h0011001110110000
`define CUBE_LUT_592 16'h0011001111111100
`define CUBE_LUT_593 16'h0011010000100100
`define CUBE_LUT_594 16'h0011010001001100
`define CUBE_LUT_595 16'h0011010001110100
`define CUBE_LUT_596 16'h0011010010011110
`define CUBE_LUT_597 16'h0011010011001000
`define CUBE_LUT_598 16'h0011010011110100
`define CUBE_LUT_599 16'h0011010100100000
`define CUBE_LUT_600 16'h0011010101001110
`define CUBE_LUT_601 16'h0011010101111100
`define CUBE_LUT_602 16'h0011010110101100
`define CUBE_LUT_603 16'h0011010111011101
`define CUBE_LUT_604 16'h0011011000001110
`define CUBE_LUT_605 16'h0011011001000001
`define CUBE_LUT_606 16'h0011011001110101
`define CUBE_LUT_607 16'h0011011010101010
`define CUBE_LUT_608 16'h0011011011100000
`define CUBE_LUT_609 16'h0011011100011000
`define CUBE_LUT_610 16'h0011011101010000
`define CUBE_LUT_611 16'h0011011110001010
`define CUBE_LUT_612 16'h0011011111000100
`define CUBE_LUT_613 16'h0011100000000000
`define CUBE_LUT_614 16'h0011100000011111
`define CUBE_LUT_615 16'h0011100000111110
`define CUBE_LUT_616 16'h0011100001011110
`define CUBE_LUT_617 16'h0011100001111110
`define CUBE_LUT_618 16'h0011100010011111
`define CUBE_LUT_619 16'h0011100011000001
`define CUBE_LUT_620 16'h0011100011100011
`define CUBE_LUT_621 16'h0011100100000110
`define CUBE_LUT_622 16'h0011100100101001
`define CUBE_LUT_623 16'h0011100101001110
`define CUBE_LUT_624 16'h0011100101110011
`define CUBE_LUT_625 16'h0011100110011000
`define CUBE_LUT_626 16'h0011100110111110
`define CUBE_LUT_627 16'h0011100111100101
`define CUBE_LUT_628 16'h0011101000001101
`define CUBE_LUT_629 16'h0011101000110101
`define CUBE_LUT_630 16'h0011101001011110
`define CUBE_LUT_631 16'h0011101010000111
`define CUBE_LUT_632 16'h0011101010110010
`define CUBE_LUT_633 16'h0011101011011101
`define CUBE_LUT_634 16'h0011101100001000
`define CUBE_LUT_635 16'h0011101100110101
`define CUBE_LUT_636 16'h0011101101100010
`define CUBE_LUT_637 16'h0011101110010000
`define CUBE_LUT_638 16'h0011101110111111
`define CUBE_LUT_639 16'h0011101111101110
`define CUBE_LUT_640 16'h0011110000001111
`define CUBE_LUT_641 16'h0011110000101000
`define CUBE_LUT_642 16'h0011110001000000
`define CUBE_LUT_643 16'h0011110001011010
`define CUBE_LUT_644 16'h0011110001110011
`define CUBE_LUT_645 16'h0011110010001101
`define CUBE_LUT_646 16'h0011110010101000
`define CUBE_LUT_647 16'h0011110011000010
`define CUBE_LUT_648 16'h0011110011011101
`define CUBE_LUT_649 16'h0011110011111001
`define CUBE_LUT_650 16'h0011110100010101
`define CUBE_LUT_651 16'h0011110100110001
`define CUBE_LUT_652 16'h0011110101001110
`define CUBE_LUT_653 16'h0011110101101011
`define CUBE_LUT_654 16'h0011110110001001
`define CUBE_LUT_655 16'h0011110110100111
`define CUBE_LUT_656 16'h0011110111000110
`define CUBE_LUT_657 16'h0011110111100100
`define CUBE_LUT_658 16'h0011111000000100
`define CUBE_LUT_659 16'h0011111000100100
`define CUBE_LUT_660 16'h0011111001000100
`define CUBE_LUT_661 16'h0011111001100100
`define CUBE_LUT_662 16'h0011111010000101
`define CUBE_LUT_663 16'h0011111010100111
`define CUBE_LUT_664 16'h0011111011001001
`define CUBE_LUT_665 16'h0011111011101011
`define CUBE_LUT_666 16'h0011111100001110
`define CUBE_LUT_667 16'h0011111100110001
`define CUBE_LUT_668 16'h0011111101010101
`define CUBE_LUT_669 16'h0011111101111001
`define CUBE_LUT_670 16'h0011111110011110
`define CUBE_LUT_671 16'h0011111111000011
`define CUBE_LUT_672 16'h0011111111101001
`define CUBE_LUT_673 16'h0100000000000111
`define CUBE_LUT_674 16'h0100000000011011
`define CUBE_LUT_675 16'h0100000000101110
`define CUBE_LUT_676 16'h0100000001000010
`define CUBE_LUT_677 16'h0100000001010110
`define CUBE_LUT_678 16'h0100000001101010
`define CUBE_LUT_679 16'h0100000001111111
`define CUBE_LUT_680 16'h0100000010010011
`define CUBE_LUT_681 16'h0100000010101000
`define CUBE_LUT_682 16'h0100000010111110
`define CUBE_LUT_683 16'h0100000011010011
`define CUBE_LUT_684 16'h0100000011101001
`define CUBE_LUT_685 16'h0100000011111111
`define CUBE_LUT_686 16'h0100000100010101
`define CUBE_LUT_687 16'h0100000100101100
`define CUBE_LUT_688 16'h0100000101000010
`define CUBE_LUT_689 16'h0100000101011001
`define CUBE_LUT_690 16'h0100000101110001
`define CUBE_LUT_691 16'h0100000110001000
`define CUBE_LUT_692 16'h0100000110100000
`define CUBE_LUT_693 16'h0100000110111000
`define CUBE_LUT_694 16'h0100000111010000
`define CUBE_LUT_695 16'h0100000111101001
`define CUBE_LUT_696 16'h0100001000000010
`define CUBE_LUT_697 16'h0100001000011011
`define CUBE_LUT_698 16'h0100001000110100
`define CUBE_LUT_699 16'h0100001001001110
`define CUBE_LUT_700 16'h0100001001101000
`define CUBE_LUT_701 16'h0100001010000010
`define CUBE_LUT_702 16'h0100001010011101
`define CUBE_LUT_703 16'h0100001010111000
`define CUBE_LUT_704 16'h0100001011010011
`define CUBE_LUT_705 16'h0100001011101110
`define CUBE_LUT_706 16'h0100001100001010
`define CUBE_LUT_707 16'h0100001100100110
`define CUBE_LUT_708 16'h0100001101000010
`define CUBE_LUT_709 16'h0100001101011110
`define CUBE_LUT_710 16'h0100001101111011
`define CUBE_LUT_711 16'h0100001110011000
`define CUBE_LUT_712 16'h0100001110110110
`define CUBE_LUT_713 16'h0100001111010011
`define CUBE_LUT_714 16'h0100001111110001
`define CUBE_LUT_715 16'h0100010000001000
`define CUBE_LUT_716 16'h0100010000010111
`define CUBE_LUT_717 16'h0100010000100110
`define CUBE_LUT_718 16'h0100010000110110
`define CUBE_LUT_719 16'h0100010001000110
`define CUBE_LUT_720 16'h0100010001010110
`define CUBE_LUT_721 16'h0100010001100110
`define CUBE_LUT_722 16'h0100010001110110
`define CUBE_LUT_723 16'h0100010010000110
`define CUBE_LUT_724 16'h0100010010010111
`define CUBE_LUT_725 16'h0100010010100111
`define CUBE_LUT_726 16'h0100010010111000
`define CUBE_LUT_727 16'h0100010011001001
`define CUBE_LUT_728 16'h0100010011011010
`define CUBE_LUT_729 16'h0100010011101100
`define CUBE_LUT_730 16'h0100010011111101
`define CUBE_LUT_731 16'h0100010100001111
`define CUBE_LUT_732 16'h0100010100100001
`define CUBE_LUT_733 16'h0100010100110010
`define CUBE_LUT_734 16'h0100010101000101
`define CUBE_LUT_735 16'h0100010101010111
`define CUBE_LUT_736 16'h0100010101101001
`define CUBE_LUT_737 16'h0100010101111100
`define CUBE_LUT_738 16'h0100010110001111
`define CUBE_LUT_739 16'h0100010110100010
`define CUBE_LUT_740 16'h0100010110110101
`define CUBE_LUT_741 16'h0100010111001000
`define CUBE_LUT_742 16'h0100010111011011
`define CUBE_LUT_743 16'h0100010111101111
`define CUBE_LUT_744 16'h0100011000000011
`define CUBE_LUT_745 16'h0100011000010111
`define CUBE_LUT_746 16'h0100011000101011
`define CUBE_LUT_747 16'h0100011000111111
`define CUBE_LUT_748 16'h0100011001010011
`define CUBE_LUT_749 16'h0100011001101000
`define CUBE_LUT_750 16'h0100011001111101
`define CUBE_LUT_751 16'h0100011010010010
`define CUBE_LUT_752 16'h0100011010100111
`define CUBE_LUT_753 16'h0100011010111100
`define CUBE_LUT_754 16'h0100011011010010
`define CUBE_LUT_755 16'h0100011011101000
`define CUBE_LUT_756 16'h0100011011111101
`define CUBE_LUT_757 16'h0100011100010011
`define CUBE_LUT_758 16'h0100011100101010
`define CUBE_LUT_759 16'h0100011101000000
`define CUBE_LUT_760 16'h0100011101010111
`define CUBE_LUT_761 16'h0100011101101101
`define CUBE_LUT_762 16'h0100011110000100
`define CUBE_LUT_763 16'h0100011110011100
`define CUBE_LUT_764 16'h0100011110110011
`define CUBE_LUT_765 16'h0100011111001010
`define CUBE_LUT_766 16'h0100011111100010
`define CUBE_LUT_767 16'h0100011111111010
`define CUBE_LUT_768 16'h0100100000001001
`define CUBE_LUT_769 16'h0100100000010101
`define CUBE_LUT_770 16'h0100100000100001
`define CUBE_LUT_771 16'h0100100000101110
`define CUBE_LUT_772 16'h0100100000111010
`define CUBE_LUT_773 16'h0100100001000111
`define CUBE_LUT_774 16'h0100100001010011
`define CUBE_LUT_775 16'h0100100001100000
`define CUBE_LUT_776 16'h0100100001101101
`define CUBE_LUT_777 16'h0100100001111010
`define CUBE_LUT_778 16'h0100100010000111
`define CUBE_LUT_779 16'h0100100010010100
`define CUBE_LUT_780 16'h0100100010100001
`define CUBE_LUT_781 16'h0100100010101110
`define CUBE_LUT_782 16'h0100100010111100
`define CUBE_LUT_783 16'h0100100011001001
`define CUBE_LUT_784 16'h0100100011010111
`define CUBE_LUT_785 16'h0100100011100100
`define CUBE_LUT_786 16'h0100100011110010
`define CUBE_LUT_787 16'h0100100100000000
`define CUBE_LUT_788 16'h0100100100001110
`define CUBE_LUT_789 16'h0100100100011100
`define CUBE_LUT_790 16'h0100100100101010
`define CUBE_LUT_791 16'h0100100100111001
`define CUBE_LUT_792 16'h0100100101000111
`define CUBE_LUT_793 16'h0100100101010101
`define CUBE_LUT_794 16'h0100100101100100
`define CUBE_LUT_795 16'h0100100101110011
`define CUBE_LUT_796 16'h0100100110000010
`define CUBE_LUT_797 16'h0100100110010001
`define CUBE_LUT_798 16'h0100100110100000
`define CUBE_LUT_799 16'h0100100110101111
`define CUBE_LUT_800 16'h0100100110111110
`define CUBE_LUT_801 16'h0100100111001101
`define CUBE_LUT_802 16'h0100100111011101
`define CUBE_LUT_803 16'h0100100111101100
`define CUBE_LUT_804 16'h0100100111111100
`define CUBE_LUT_805 16'h0100101000001100
`define CUBE_LUT_806 16'h0100101000011100
`define CUBE_LUT_807 16'h0100101000101100
`define CUBE_LUT_808 16'h0100101000111100
`define CUBE_LUT_809 16'h0100101001001100
`define CUBE_LUT_810 16'h0100101001011100
`define CUBE_LUT_811 16'h0100101001101101
`define CUBE_LUT_812 16'h0100101001111101
`define CUBE_LUT_813 16'h0100101010001110
`define CUBE_LUT_814 16'h0100101010011110
`define CUBE_LUT_815 16'h0100101010101111
`define CUBE_LUT_816 16'h0100101011000000
`define CUBE_LUT_817 16'h0100101011010001
`define CUBE_LUT_818 16'h0100101011100011
`define CUBE_LUT_819 16'h0100101011110100
`define CUBE_LUT_820 16'h0100101100000101
`define CUBE_LUT_821 16'h0100101100010111
`define CUBE_LUT_822 16'h0100101100101000
`define CUBE_LUT_823 16'h0100101100111010
`define CUBE_LUT_824 16'h0100101101001100
`define CUBE_LUT_825 16'h0100101101011110
`define CUBE_LUT_826 16'h0100101101110000
`define CUBE_LUT_827 16'h0100101110000010
`define CUBE_LUT_828 16'h0100101110010101
`define CUBE_LUT_829 16'h0100101110100111
`define CUBE_LUT_830 16'h0100101110111010
`define CUBE_LUT_831 16'h0100101111001100
`define CUBE_LUT_832 16'h0100101111011111
`define CUBE_LUT_833 16'h0100101111110010
`define CUBE_LUT_834 16'h0100110000000011
`define CUBE_LUT_835 16'h0100110000001100
`define CUBE_LUT_836 16'h0100110000010110
`define CUBE_LUT_837 16'h0100110000100000
`define CUBE_LUT_838 16'h0100110000101001
`define CUBE_LUT_839 16'h0100110000110011
`define CUBE_LUT_840 16'h0100110000111101
`define CUBE_LUT_841 16'h0100110001000111
`define CUBE_LUT_842 16'h0100110001010001
`define CUBE_LUT_843 16'h0100110001011011
`define CUBE_LUT_844 16'h0100110001100101
`define CUBE_LUT_845 16'h0100110001101111
`define CUBE_LUT_846 16'h0100110001111010
`define CUBE_LUT_847 16'h0100110010000100
`define CUBE_LUT_848 16'h0100110010001110
`define CUBE_LUT_849 16'h0100110010011001
`define CUBE_LUT_850 16'h0100110010100011
`define CUBE_LUT_851 16'h0100110010101110
`define CUBE_LUT_852 16'h0100110010111000
`define CUBE_LUT_853 16'h0100110011000011
`define CUBE_LUT_854 16'h0100110011001110
`define CUBE_LUT_855 16'h0100110011011001
`define CUBE_LUT_856 16'h0100110011100011
`define CUBE_LUT_857 16'h0100110011101110
`define CUBE_LUT_858 16'h0100110011111001
`define CUBE_LUT_859 16'h0100110100000100
`define CUBE_LUT_860 16'h0100110100001111
`define CUBE_LUT_861 16'h0100110100011011
`define CUBE_LUT_862 16'h0100110100100110
`define CUBE_LUT_863 16'h0100110100110001
`define CUBE_LUT_864 16'h0100110100111101
`define CUBE_LUT_865 16'h0100110101001000
`define CUBE_LUT_866 16'h0100110101010100
`define CUBE_LUT_867 16'h0100110101011111
`define CUBE_LUT_868 16'h0100110101101011
`define CUBE_LUT_869 16'h0100110101110110
`define CUBE_LUT_870 16'h0100110110000010
`define CUBE_LUT_871 16'h0100110110001110
`define CUBE_LUT_872 16'h0100110110011010
`define CUBE_LUT_873 16'h0100110110100110
`define CUBE_LUT_874 16'h0100110110110010
`define CUBE_LUT_875 16'h0100110110111110
`define CUBE_LUT_876 16'h0100110111001010
`define CUBE_LUT_877 16'h0100110111010110
`define CUBE_LUT_878 16'h0100110111100011
`define CUBE_LUT_879 16'h0100110111101111
`define CUBE_LUT_880 16'h0100110111111100
`define CUBE_LUT_881 16'h0100111000001000
`define CUBE_LUT_882 16'h0100111000010101
`define CUBE_LUT_883 16'h0100111000100001
`define CUBE_LUT_884 16'h0100111000101110
`define CUBE_LUT_885 16'h0100111000111011
`define CUBE_LUT_886 16'h0100111001001000
`define CUBE_LUT_887 16'h0100111001010101
`define CUBE_LUT_888 16'h0100111001100001
`define CUBE_LUT_889 16'h0100111001101111
`define CUBE_LUT_890 16'h0100111001111100
`define CUBE_LUT_891 16'h0100111010001001
`define CUBE_LUT_892 16'h0100111010010110
`define CUBE_LUT_893 16'h0100111010100011
`define CUBE_LUT_894 16'h0100111010110001
`define CUBE_LUT_895 16'h0100111010111110
`define CUBE_LUT_896 16'h0100111011001100
`define CUBE_LUT_897 16'h0100111011011001
`define CUBE_LUT_898 16'h0100111011100111
`define CUBE_LUT_899 16'h0100111011110101
`define CUBE_LUT_900 16'h0100111100000011
`define CUBE_LUT_901 16'h0100111100010001
`define CUBE_LUT_902 16'h0100111100011111
`define CUBE_LUT_903 16'h0100111100101101
`define CUBE_LUT_904 16'h0100111100111011
`define CUBE_LUT_905 16'h0100111101001001
`define CUBE_LUT_906 16'h0100111101010111
`define CUBE_LUT_907 16'h0100111101100101
`define CUBE_LUT_908 16'h0100111101110100
`define CUBE_LUT_909 16'h0100111110000010
`define CUBE_LUT_910 16'h0100111110010001
`define CUBE_LUT_911 16'h0100111110100000
`define CUBE_LUT_912 16'h0100111110101110
`define CUBE_LUT_913 16'h0100111110111101
`define CUBE_LUT_914 16'h0100111111001100
`define CUBE_LUT_915 16'h0100111111011011
`define CUBE_LUT_916 16'h0100111111101010
`define CUBE_LUT_917 16'h0100111111111001
`define CUBE_LUT_918 16'h0101000000000100
`define CUBE_LUT_919 16'h0101000000001100
`define CUBE_LUT_920 16'h0101000000010011
`define CUBE_LUT_921 16'h0101000000011011
`define CUBE_LUT_922 16'h0101000000100011
`define CUBE_LUT_923 16'h0101000000101010
`define CUBE_LUT_924 16'h0101000000110010
`define CUBE_LUT_925 16'h0101000000111010
`define CUBE_LUT_926 16'h0101000001000010
`define CUBE_LUT_927 16'h0101000001001010
`define CUBE_LUT_928 16'h0101000001010010
`define CUBE_LUT_929 16'h0101000001011010
`define CUBE_LUT_930 16'h0101000001100010
`define CUBE_LUT_931 16'h0101000001101010
`define CUBE_LUT_932 16'h0101000001110010
`define CUBE_LUT_933 16'h0101000001111010
`define CUBE_LUT_934 16'h0101000010000010
`define CUBE_LUT_935 16'h0101000010001010
`define CUBE_LUT_936 16'h0101000010010011
`define CUBE_LUT_937 16'h0101000010011011
`define CUBE_LUT_938 16'h0101000010100011
`define CUBE_LUT_939 16'h0101000010101100
`define CUBE_LUT_940 16'h0101000010110100
`define CUBE_LUT_941 16'h0101000010111101
`define CUBE_LUT_942 16'h0101000011000101
`define CUBE_LUT_943 16'h0101000011001110
`define CUBE_LUT_944 16'h0101000011010110
`define CUBE_LUT_945 16'h0101000011011111
`define CUBE_LUT_946 16'h0101000011100111
`define CUBE_LUT_947 16'h0101000011110000
`define CUBE_LUT_948 16'h0101000011111001
`define CUBE_LUT_949 16'h0101000100000010
`define CUBE_LUT_950 16'h0101000100001010
`define CUBE_LUT_951 16'h0101000100010011
`define CUBE_LUT_952 16'h0101000100011100
`define CUBE_LUT_953 16'h0101000100100101
`define CUBE_LUT_954 16'h0101000100101110
`define CUBE_LUT_955 16'h0101000100110111
`define CUBE_LUT_956 16'h0101000101000000
`define CUBE_LUT_957 16'h0101000101001001
`define CUBE_LUT_958 16'h0101000101010010
`define CUBE_LUT_959 16'h0101000101011011
`define CUBE_LUT_960 16'h0101000101100101
`define CUBE_LUT_961 16'h0101000101101110
`define CUBE_LUT_962 16'h0101000101110111
`define CUBE_LUT_963 16'h0101000110000001
`define CUBE_LUT_964 16'h0101000110001010
`define CUBE_LUT_965 16'h0101000110010011
`define CUBE_LUT_966 16'h0101000110011101
`define CUBE_LUT_967 16'h0101000110100110
`define CUBE_LUT_968 16'h0101000110110000
`define CUBE_LUT_969 16'h0101000110111001
`define CUBE_LUT_970 16'h0101000111000011
`define CUBE_LUT_971 16'h0101000111001101
`define CUBE_LUT_972 16'h0101000111010110
`define CUBE_LUT_973 16'h0101000111100000
`define CUBE_LUT_974 16'h0101000111101010
`define CUBE_LUT_975 16'h0101000111110100
`define CUBE_LUT_976 16'h0101000111111110
`define CUBE_LUT_977 16'h0101001000001000
`define CUBE_LUT_978 16'h0101001000010010
`define CUBE_LUT_979 16'h0101001000011100
`define CUBE_LUT_980 16'h0101001000100110
`define CUBE_LUT_981 16'h0101001000110000
`define CUBE_LUT_982 16'h0101001000111010
`define CUBE_LUT_983 16'h0101001001000100
`define CUBE_LUT_984 16'h0101001001001110
`define CUBE_LUT_985 16'h0101001001011001
`define CUBE_LUT_986 16'h0101001001100011
`define CUBE_LUT_987 16'h0101001001101101
`define CUBE_LUT_988 16'h0101001001111000
`define CUBE_LUT_989 16'h0101001010000010
`define CUBE_LUT_990 16'h0101001010001101
`define CUBE_LUT_991 16'h0101001010010111
`define CUBE_LUT_992 16'h0101001010100010
`define CUBE_LUT_993 16'h0101001010101100
`define CUBE_LUT_994 16'h0101001010110111
`define CUBE_LUT_995 16'h0101001011000010
`define CUBE_LUT_996 16'h0101001011001101
`define CUBE_LUT_997 16'h0101001011010111
`define CUBE_LUT_998 16'h0101001011100010
`define CUBE_LUT_999 16'h0101001011101101
`define CUBE_LUT_1000 16'h0101001011111000
`define CUBE_LUT_1001 16'h0101001100000011
`define CUBE_LUT_1002 16'h0101001100001110
`define CUBE_LUT_1003 16'h0101001100011001
`define CUBE_LUT_1004 16'h0101001100100100
`define CUBE_LUT_1005 16'h0101001100101111
`define CUBE_LUT_1006 16'h0101001100111011
`define CUBE_LUT_1007 16'h0101001101000110
`define CUBE_LUT_1008 16'h0101001101010001
`define CUBE_LUT_1009 16'h0101001101011100
`define CUBE_LUT_1010 16'h0101001101101000
`define CUBE_LUT_1011 16'h0101001101110011
`define CUBE_LUT_1012 16'h0101001101111111
`define CUBE_LUT_1013 16'h0101001110001010
`define CUBE_LUT_1014 16'h0101001110010110
`define CUBE_LUT_1015 16'h0101001110100001
`define CUBE_LUT_1016 16'h0101001110101101
`define CUBE_LUT_1017 16'h0101001110111001
`define CUBE_LUT_1018 16'h0101001111000101
`define CUBE_LUT_1019 16'h0101001111010000
`define CUBE_LUT_1020 16'h0101001111011100
`define CUBE_LUT_1021 16'h0101001111101000
`define CUBE_LUT_1022 16'h0101001111110100
`define CUBE_LUT_1023 16'h0101010000000000
