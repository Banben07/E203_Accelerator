`define TANH_LUT_SIZE 4280
`define TANH_LUT_BITS 13
`define TANH_LUT_0000 16'h0000
`define TANH_LUT_0008 16'h0008
`define TANH_LUT_0010 16'h0010
`define TANH_LUT_0018 16'h0018
`define TANH_LUT_0020 16'h0020
`define TANH_LUT_0028 16'h0028
`define TANH_LUT_0030 16'h0030
`define TANH_LUT_0038 16'h0038
`define TANH_LUT_0040 16'h0040
`define TANH_LUT_0048 16'h0048
`define TANH_LUT_0050 16'h0050
`define TANH_LUT_0058 16'h0058
`define TANH_LUT_0060 16'h0060
`define TANH_LUT_0068 16'h0068
`define TANH_LUT_0070 16'h0070
`define TANH_LUT_0078 16'h0078
`define TANH_LUT_0080 16'h0080
`define TANH_LUT_0088 16'h0088
`define TANH_LUT_0090 16'h0090
`define TANH_LUT_0098 16'h0098
`define TANH_LUT_00A0 16'h00A0
`define TANH_LUT_00A8 16'h00A8
`define TANH_LUT_00B0 16'h00B0
`define TANH_LUT_00B8 16'h00B8
`define TANH_LUT_00C0 16'h00C0
`define TANH_LUT_00C8 16'h00C8
`define TANH_LUT_00D0 16'h00D0
`define TANH_LUT_00D8 16'h00D8
`define TANH_LUT_00E0 16'h00E0
`define TANH_LUT_00E8 16'h00E8
`define TANH_LUT_00F0 16'h00F0
`define TANH_LUT_00F8 16'h00F8
`define TANH_LUT_0100 16'h0100
`define TANH_LUT_0108 16'h0108
`define TANH_LUT_0110 16'h0110
`define TANH_LUT_0118 16'h0118
`define TANH_LUT_0120 16'h0120
`define TANH_LUT_0128 16'h0128
`define TANH_LUT_0130 16'h0130
`define TANH_LUT_0138 16'h0138
`define TANH_LUT_0140 16'h0140
`define TANH_LUT_0148 16'h0148
`define TANH_LUT_0150 16'h0150
`define TANH_LUT_0158 16'h0158
`define TANH_LUT_0160 16'h0160
`define TANH_LUT_0168 16'h0168
`define TANH_LUT_0170 16'h0170
`define TANH_LUT_0178 16'h0178
`define TANH_LUT_0180 16'h0180
`define TANH_LUT_0188 16'h0188
`define TANH_LUT_0190 16'h0190
`define TANH_LUT_0198 16'h0198
`define TANH_LUT_01A0 16'h01A0
`define TANH_LUT_01A8 16'h01A8
`define TANH_LUT_01B0 16'h01B0
`define TANH_LUT_01B8 16'h01B8
`define TANH_LUT_01C0 16'h01C0
`define TANH_LUT_01C8 16'h01C8
`define TANH_LUT_01D0 16'h01D0
`define TANH_LUT_01D8 16'h01D8
`define TANH_LUT_01E0 16'h01E0
`define TANH_LUT_01E8 16'h01E8
`define TANH_LUT_01F0 16'h01F0
`define TANH_LUT_01F8 16'h01F8
`define TANH_LUT_0200 16'h0200
`define TANH_LUT_0208 16'h0208
`define TANH_LUT_0210 16'h0210
`define TANH_LUT_0218 16'h0218
`define TANH_LUT_0220 16'h0220
`define TANH_LUT_0228 16'h0228
`define TANH_LUT_0230 16'h0230
`define TANH_LUT_0238 16'h0238
`define TANH_LUT_0240 16'h0240
`define TANH_LUT_0248 16'h0248
`define TANH_LUT_0250 16'h0250
`define TANH_LUT_0258 16'h0258
`define TANH_LUT_0260 16'h0260
`define TANH_LUT_0268 16'h0268
`define TANH_LUT_0270 16'h0270
`define TANH_LUT_0278 16'h0278
`define TANH_LUT_0280 16'h0280
`define TANH_LUT_0288 16'h0288
`define TANH_LUT_0290 16'h0290
`define TANH_LUT_0298 16'h0298
`define TANH_LUT_02A0 16'h02A0
`define TANH_LUT_02A8 16'h02A8
`define TANH_LUT_02B0 16'h02B0
`define TANH_LUT_02B8 16'h02B8
`define TANH_LUT_02C0 16'h02C0
`define TANH_LUT_02C8 16'h02C8
`define TANH_LUT_02D0 16'h02D0
`define TANH_LUT_02D8 16'h02D8
`define TANH_LUT_02E0 16'h02E0
`define TANH_LUT_02E8 16'h02E8
`define TANH_LUT_02F0 16'h02F0
`define TANH_LUT_02F8 16'h02F8
`define TANH_LUT_0300 16'h0300
`define TANH_LUT_0308 16'h0308
`define TANH_LUT_0310 16'h0310
`define TANH_LUT_0318 16'h0318
`define TANH_LUT_0320 16'h0320
`define TANH_LUT_0328 16'h0328
`define TANH_LUT_0330 16'h0330
`define TANH_LUT_0338 16'h0338
`define TANH_LUT_0340 16'h0340
`define TANH_LUT_0348 16'h0348
`define TANH_LUT_0350 16'h0350
`define TANH_LUT_0358 16'h0358
`define TANH_LUT_0360 16'h0360
`define TANH_LUT_0368 16'h0368
`define TANH_LUT_0370 16'h0370
`define TANH_LUT_0378 16'h0378
`define TANH_LUT_0380 16'h0380
`define TANH_LUT_0388 16'h0388
`define TANH_LUT_0390 16'h0390
`define TANH_LUT_0398 16'h0398
`define TANH_LUT_03A0 16'h03A0
`define TANH_LUT_03A8 16'h03A8
`define TANH_LUT_03B0 16'h03B0
`define TANH_LUT_03B8 16'h03B8
`define TANH_LUT_03C0 16'h03C0
`define TANH_LUT_03C8 16'h03C8
`define TANH_LUT_03D0 16'h03D0
`define TANH_LUT_03D8 16'h03D8
`define TANH_LUT_03E0 16'h03E0
`define TANH_LUT_03E8 16'h03E8
`define TANH_LUT_03F0 16'h03F0
`define TANH_LUT_03F8 16'h03F8
`define TANH_LUT_0400 16'h0400
`define TANH_LUT_0408 16'h0408
`define TANH_LUT_0410 16'h0410
`define TANH_LUT_0418 16'h0418
`define TANH_LUT_0420 16'h0420
`define TANH_LUT_0428 16'h0428
`define TANH_LUT_0430 16'h0430
`define TANH_LUT_0438 16'h0438
`define TANH_LUT_0440 16'h0440
`define TANH_LUT_0448 16'h0448
`define TANH_LUT_0450 16'h0450
`define TANH_LUT_0458 16'h0458
`define TANH_LUT_0460 16'h0460
`define TANH_LUT_0468 16'h0468
`define TANH_LUT_0470 16'h0470
`define TANH_LUT_0478 16'h0478
`define TANH_LUT_0480 16'h0480
`define TANH_LUT_0488 16'h0488
`define TANH_LUT_0490 16'h0490
`define TANH_LUT_0498 16'h0498
`define TANH_LUT_04A0 16'h04A0
`define TANH_LUT_04A8 16'h04A8
`define TANH_LUT_04B0 16'h04B0
`define TANH_LUT_04B8 16'h04B8
`define TANH_LUT_04C0 16'h04C0
`define TANH_LUT_04C8 16'h04C8
`define TANH_LUT_04D0 16'h04D0
`define TANH_LUT_04D8 16'h04D8
`define TANH_LUT_04E0 16'h04E0
`define TANH_LUT_04E8 16'h04E8
`define TANH_LUT_04F0 16'h04F0
`define TANH_LUT_04F8 16'h04F8
`define TANH_LUT_0500 16'h0500
`define TANH_LUT_0508 16'h0508
`define TANH_LUT_0510 16'h0510
`define TANH_LUT_0518 16'h0518
`define TANH_LUT_0520 16'h0520
`define TANH_LUT_0528 16'h0528
`define TANH_LUT_0530 16'h0530
`define TANH_LUT_0538 16'h0538
`define TANH_LUT_0540 16'h0540
`define TANH_LUT_0548 16'h0548
`define TANH_LUT_0550 16'h0550
`define TANH_LUT_0558 16'h0558
`define TANH_LUT_0560 16'h0560
`define TANH_LUT_0568 16'h0568
`define TANH_LUT_0570 16'h0570
`define TANH_LUT_0578 16'h0578
`define TANH_LUT_0580 16'h0580
`define TANH_LUT_0588 16'h0588
`define TANH_LUT_0590 16'h0590
`define TANH_LUT_0598 16'h0598
`define TANH_LUT_05A0 16'h05A0
`define TANH_LUT_05A8 16'h05A8
`define TANH_LUT_05B0 16'h05B0
`define TANH_LUT_05B8 16'h05B8
`define TANH_LUT_05C0 16'h05C0
`define TANH_LUT_05C8 16'h05C8
`define TANH_LUT_05D0 16'h05D0
`define TANH_LUT_05D8 16'h05D8
`define TANH_LUT_05E0 16'h05E0
`define TANH_LUT_05E8 16'h05E8
`define TANH_LUT_05F0 16'h05F0
`define TANH_LUT_05F8 16'h05F8
`define TANH_LUT_0600 16'h0600
`define TANH_LUT_0608 16'h0608
`define TANH_LUT_0610 16'h0610
`define TANH_LUT_0618 16'h0618
`define TANH_LUT_0620 16'h0620
`define TANH_LUT_0628 16'h0628
`define TANH_LUT_0630 16'h0630
`define TANH_LUT_0638 16'h0638
`define TANH_LUT_0640 16'h0640
`define TANH_LUT_0648 16'h0648
`define TANH_LUT_0650 16'h0650
`define TANH_LUT_0658 16'h0658
`define TANH_LUT_0660 16'h0660
`define TANH_LUT_0668 16'h0668
`define TANH_LUT_0670 16'h0670
`define TANH_LUT_0678 16'h0678
`define TANH_LUT_0680 16'h0680
`define TANH_LUT_0688 16'h0688
`define TANH_LUT_0690 16'h0690
`define TANH_LUT_0698 16'h0698
`define TANH_LUT_06A0 16'h06A0
`define TANH_LUT_06A8 16'h06A8
`define TANH_LUT_06B0 16'h06B0
`define TANH_LUT_06B8 16'h06B8
`define TANH_LUT_06C0 16'h06C0
`define TANH_LUT_06C8 16'h06C8
`define TANH_LUT_06D0 16'h06D0
`define TANH_LUT_06D8 16'h06D8
`define TANH_LUT_06E0 16'h06E0
`define TANH_LUT_06E8 16'h06E8
`define TANH_LUT_06F0 16'h06F0
`define TANH_LUT_06F8 16'h06F8
`define TANH_LUT_0700 16'h0700
`define TANH_LUT_0708 16'h0708
`define TANH_LUT_0710 16'h0710
`define TANH_LUT_0718 16'h0718
`define TANH_LUT_0720 16'h0720
`define TANH_LUT_0728 16'h0728
`define TANH_LUT_0730 16'h0730
`define TANH_LUT_0738 16'h0738
`define TANH_LUT_0740 16'h0740
`define TANH_LUT_0748 16'h0748
`define TANH_LUT_0750 16'h0750
`define TANH_LUT_0758 16'h0758
`define TANH_LUT_0760 16'h0760
`define TANH_LUT_0768 16'h0768
`define TANH_LUT_0770 16'h0770
`define TANH_LUT_0778 16'h0778
`define TANH_LUT_0780 16'h0780
`define TANH_LUT_0788 16'h0788
`define TANH_LUT_0790 16'h0790
`define TANH_LUT_0798 16'h0798
`define TANH_LUT_07A0 16'h07A0
`define TANH_LUT_07A8 16'h07A8
`define TANH_LUT_07B0 16'h07B0
`define TANH_LUT_07B8 16'h07B8
`define TANH_LUT_07C0 16'h07C0
`define TANH_LUT_07C8 16'h07C8
`define TANH_LUT_07D0 16'h07D0
`define TANH_LUT_07D8 16'h07D8
`define TANH_LUT_07E0 16'h07E0
`define TANH_LUT_07E8 16'h07E8
`define TANH_LUT_07F0 16'h07F0
`define TANH_LUT_07F8 16'h07F8
`define TANH_LUT_0800 16'h0800
`define TANH_LUT_0808 16'h0808
`define TANH_LUT_0810 16'h0810
`define TANH_LUT_0818 16'h0818
`define TANH_LUT_0820 16'h0820
`define TANH_LUT_0828 16'h0828
`define TANH_LUT_0830 16'h0830
`define TANH_LUT_0838 16'h0838
`define TANH_LUT_0840 16'h0840
`define TANH_LUT_0848 16'h0848
`define TANH_LUT_0850 16'h0850
`define TANH_LUT_0858 16'h0858
`define TANH_LUT_0860 16'h0860
`define TANH_LUT_0868 16'h0868
`define TANH_LUT_0870 16'h0870
`define TANH_LUT_0878 16'h0878
`define TANH_LUT_0880 16'h0880
`define TANH_LUT_0888 16'h0888
`define TANH_LUT_0890 16'h0890
`define TANH_LUT_0898 16'h0898
`define TANH_LUT_08A0 16'h08A0
`define TANH_LUT_08A8 16'h08A8
`define TANH_LUT_08B0 16'h08B0
`define TANH_LUT_08B8 16'h08B8
`define TANH_LUT_08C0 16'h08C0
`define TANH_LUT_08C8 16'h08C8
`define TANH_LUT_08D0 16'h08D0
`define TANH_LUT_08D8 16'h08D8
`define TANH_LUT_08E0 16'h08E0
`define TANH_LUT_08E8 16'h08E8
`define TANH_LUT_08F0 16'h08F0
`define TANH_LUT_08F8 16'h08F8
`define TANH_LUT_0900 16'h0900
`define TANH_LUT_0908 16'h0908
`define TANH_LUT_0910 16'h0910
`define TANH_LUT_0918 16'h0918
`define TANH_LUT_0920 16'h0920
`define TANH_LUT_0928 16'h0928
`define TANH_LUT_0930 16'h0930
`define TANH_LUT_0938 16'h0938
`define TANH_LUT_0940 16'h0940
`define TANH_LUT_0948 16'h0948
`define TANH_LUT_0950 16'h0950
`define TANH_LUT_0958 16'h0958
`define TANH_LUT_0960 16'h0960
`define TANH_LUT_0968 16'h0968
`define TANH_LUT_0970 16'h0970
`define TANH_LUT_0978 16'h0978
`define TANH_LUT_0980 16'h0980
`define TANH_LUT_0988 16'h0988
`define TANH_LUT_0990 16'h0990
`define TANH_LUT_0998 16'h0998
`define TANH_LUT_09A0 16'h09A0
`define TANH_LUT_09A8 16'h09A8
`define TANH_LUT_09B0 16'h09B0
`define TANH_LUT_09B8 16'h09B8
`define TANH_LUT_09C0 16'h09C0
`define TANH_LUT_09C8 16'h09C8
`define TANH_LUT_09D0 16'h09D0
`define TANH_LUT_09D8 16'h09D8
`define TANH_LUT_09E0 16'h09E0
`define TANH_LUT_09E8 16'h09E8
`define TANH_LUT_09F0 16'h09F0
`define TANH_LUT_09F8 16'h09F8
`define TANH_LUT_0A00 16'h0A00
`define TANH_LUT_0A08 16'h0A08
`define TANH_LUT_0A10 16'h0A10
`define TANH_LUT_0A18 16'h0A18
`define TANH_LUT_0A20 16'h0A20
`define TANH_LUT_0A28 16'h0A28
`define TANH_LUT_0A30 16'h0A30
`define TANH_LUT_0A38 16'h0A38
`define TANH_LUT_0A40 16'h0A40
`define TANH_LUT_0A48 16'h0A48
`define TANH_LUT_0A50 16'h0A50
`define TANH_LUT_0A58 16'h0A58
`define TANH_LUT_0A60 16'h0A60
`define TANH_LUT_0A68 16'h0A68
`define TANH_LUT_0A70 16'h0A70
`define TANH_LUT_0A78 16'h0A78
`define TANH_LUT_0A80 16'h0A80
`define TANH_LUT_0A88 16'h0A88
`define TANH_LUT_0A90 16'h0A90
`define TANH_LUT_0A98 16'h0A98
`define TANH_LUT_0AA0 16'h0AA0
`define TANH_LUT_0AA8 16'h0AA8
`define TANH_LUT_0AB0 16'h0AB0
`define TANH_LUT_0AB8 16'h0AB8
`define TANH_LUT_0AC0 16'h0AC0
`define TANH_LUT_0AC8 16'h0AC8
`define TANH_LUT_0AD0 16'h0AD0
`define TANH_LUT_0AD8 16'h0AD8
`define TANH_LUT_0AE0 16'h0AE0
`define TANH_LUT_0AE8 16'h0AE8
`define TANH_LUT_0AF0 16'h0AF0
`define TANH_LUT_0AF8 16'h0AF8
`define TANH_LUT_0B00 16'h0B00
`define TANH_LUT_0B08 16'h0B08
`define TANH_LUT_0B10 16'h0B10
`define TANH_LUT_0B18 16'h0B18
`define TANH_LUT_0B20 16'h0B20
`define TANH_LUT_0B28 16'h0B28
`define TANH_LUT_0B30 16'h0B30
`define TANH_LUT_0B38 16'h0B38
`define TANH_LUT_0B40 16'h0B40
`define TANH_LUT_0B48 16'h0B48
`define TANH_LUT_0B50 16'h0B50
`define TANH_LUT_0B58 16'h0B58
`define TANH_LUT_0B60 16'h0B60
`define TANH_LUT_0B68 16'h0B68
`define TANH_LUT_0B70 16'h0B70
`define TANH_LUT_0B78 16'h0B78
`define TANH_LUT_0B80 16'h0B80
`define TANH_LUT_0B88 16'h0B88
`define TANH_LUT_0B90 16'h0B90
`define TANH_LUT_0B98 16'h0B98
`define TANH_LUT_0BA0 16'h0BA0
`define TANH_LUT_0BA8 16'h0BA8
`define TANH_LUT_0BB0 16'h0BB0
`define TANH_LUT_0BB8 16'h0BB8
`define TANH_LUT_0BC0 16'h0BC0
`define TANH_LUT_0BC8 16'h0BC8
`define TANH_LUT_0BD0 16'h0BD0
`define TANH_LUT_0BD8 16'h0BD8
`define TANH_LUT_0BE0 16'h0BE0
`define TANH_LUT_0BE8 16'h0BE8
`define TANH_LUT_0BF0 16'h0BF0
`define TANH_LUT_0BF8 16'h0BF8
`define TANH_LUT_0C00 16'h0C00
`define TANH_LUT_0C08 16'h0C08
`define TANH_LUT_0C10 16'h0C10
`define TANH_LUT_0C18 16'h0C18
`define TANH_LUT_0C20 16'h0C20
`define TANH_LUT_0C28 16'h0C28
`define TANH_LUT_0C30 16'h0C30
`define TANH_LUT_0C38 16'h0C38
`define TANH_LUT_0C40 16'h0C40
`define TANH_LUT_0C48 16'h0C48
`define TANH_LUT_0C50 16'h0C50
`define TANH_LUT_0C58 16'h0C58
`define TANH_LUT_0C60 16'h0C60
`define TANH_LUT_0C68 16'h0C68
`define TANH_LUT_0C70 16'h0C70
`define TANH_LUT_0C78 16'h0C78
`define TANH_LUT_0C80 16'h0C80
`define TANH_LUT_0C88 16'h0C88
`define TANH_LUT_0C90 16'h0C90
`define TANH_LUT_0C98 16'h0C98
`define TANH_LUT_0CA0 16'h0CA0
`define TANH_LUT_0CA8 16'h0CA8
`define TANH_LUT_0CB0 16'h0CB0
`define TANH_LUT_0CB8 16'h0CB8
`define TANH_LUT_0CC0 16'h0CC0
`define TANH_LUT_0CC8 16'h0CC8
`define TANH_LUT_0CD0 16'h0CD0
`define TANH_LUT_0CD8 16'h0CD8
`define TANH_LUT_0CE0 16'h0CE0
`define TANH_LUT_0CE8 16'h0CE8
`define TANH_LUT_0CF0 16'h0CF0
`define TANH_LUT_0CF8 16'h0CF8
`define TANH_LUT_0D00 16'h0D00
`define TANH_LUT_0D08 16'h0D08
`define TANH_LUT_0D10 16'h0D10
`define TANH_LUT_0D18 16'h0D18
`define TANH_LUT_0D20 16'h0D20
`define TANH_LUT_0D28 16'h0D28
`define TANH_LUT_0D30 16'h0D30
`define TANH_LUT_0D38 16'h0D38
`define TANH_LUT_0D40 16'h0D40
`define TANH_LUT_0D48 16'h0D48
`define TANH_LUT_0D50 16'h0D50
`define TANH_LUT_0D58 16'h0D58
`define TANH_LUT_0D60 16'h0D60
`define TANH_LUT_0D68 16'h0D68
`define TANH_LUT_0D70 16'h0D70
`define TANH_LUT_0D78 16'h0D78
`define TANH_LUT_0D80 16'h0D80
`define TANH_LUT_0D88 16'h0D88
`define TANH_LUT_0D90 16'h0D90
`define TANH_LUT_0D98 16'h0D98
`define TANH_LUT_0DA0 16'h0DA0
`define TANH_LUT_0DA8 16'h0DA8
`define TANH_LUT_0DB0 16'h0DB0
`define TANH_LUT_0DB8 16'h0DB8
`define TANH_LUT_0DC0 16'h0DC0
`define TANH_LUT_0DC8 16'h0DC8
`define TANH_LUT_0DD0 16'h0DD0
`define TANH_LUT_0DD8 16'h0DD8
`define TANH_LUT_0DE0 16'h0DE0
`define TANH_LUT_0DE8 16'h0DE8
`define TANH_LUT_0DF0 16'h0DF0
`define TANH_LUT_0DF8 16'h0DF8
`define TANH_LUT_0E00 16'h0E00
`define TANH_LUT_0E08 16'h0E08
`define TANH_LUT_0E10 16'h0E10
`define TANH_LUT_0E18 16'h0E18
`define TANH_LUT_0E20 16'h0E20
`define TANH_LUT_0E28 16'h0E28
`define TANH_LUT_0E30 16'h0E30
`define TANH_LUT_0E38 16'h0E38
`define TANH_LUT_0E40 16'h0E40
`define TANH_LUT_0E48 16'h0E48
`define TANH_LUT_0E50 16'h0E50
`define TANH_LUT_0E58 16'h0E58
`define TANH_LUT_0E60 16'h0E60
`define TANH_LUT_0E68 16'h0E68
`define TANH_LUT_0E70 16'h0E70
`define TANH_LUT_0E78 16'h0E78
`define TANH_LUT_0E80 16'h0E80
`define TANH_LUT_0E88 16'h0E88
`define TANH_LUT_0E90 16'h0E90
`define TANH_LUT_0E98 16'h0E98
`define TANH_LUT_0EA0 16'h0EA0
`define TANH_LUT_0EA8 16'h0EA8
`define TANH_LUT_0EB0 16'h0EB0
`define TANH_LUT_0EB8 16'h0EB8
`define TANH_LUT_0EC0 16'h0EC0
`define TANH_LUT_0EC8 16'h0EC8
`define TANH_LUT_0ED0 16'h0ED0
`define TANH_LUT_0ED8 16'h0ED8
`define TANH_LUT_0EE0 16'h0EE0
`define TANH_LUT_0EE8 16'h0EE8
`define TANH_LUT_0EF0 16'h0EF0
`define TANH_LUT_0EF8 16'h0EF8
`define TANH_LUT_0F00 16'h0F00
`define TANH_LUT_0F08 16'h0F08
`define TANH_LUT_0F10 16'h0F10
`define TANH_LUT_0F18 16'h0F18
`define TANH_LUT_0F20 16'h0F20
`define TANH_LUT_0F28 16'h0F28
`define TANH_LUT_0F30 16'h0F30
`define TANH_LUT_0F38 16'h0F38
`define TANH_LUT_0F40 16'h0F40
`define TANH_LUT_0F48 16'h0F48
`define TANH_LUT_0F50 16'h0F50
`define TANH_LUT_0F58 16'h0F58
`define TANH_LUT_0F60 16'h0F60
`define TANH_LUT_0F68 16'h0F68
`define TANH_LUT_0F70 16'h0F70
`define TANH_LUT_0F78 16'h0F78
`define TANH_LUT_0F80 16'h0F80
`define TANH_LUT_0F88 16'h0F88
`define TANH_LUT_0F90 16'h0F90
`define TANH_LUT_0F98 16'h0F98
`define TANH_LUT_0FA0 16'h0FA0
`define TANH_LUT_0FA8 16'h0FA8
`define TANH_LUT_0FB0 16'h0FB0
`define TANH_LUT_0FB8 16'h0FB8
`define TANH_LUT_0FC0 16'h0FC0
`define TANH_LUT_0FC8 16'h0FC8
`define TANH_LUT_0FD0 16'h0FD0
`define TANH_LUT_0FD8 16'h0FD8
`define TANH_LUT_0FE0 16'h0FE0
`define TANH_LUT_0FE8 16'h0FE8
`define TANH_LUT_0FF0 16'h0FF0
`define TANH_LUT_0FF8 16'h0FF8
`define TANH_LUT_1000 16'h1000
`define TANH_LUT_1008 16'h1008
`define TANH_LUT_1010 16'h1010
`define TANH_LUT_1018 16'h1018
`define TANH_LUT_1020 16'h1020
`define TANH_LUT_1028 16'h1028
`define TANH_LUT_1030 16'h1030
`define TANH_LUT_1038 16'h1038
`define TANH_LUT_1040 16'h1040
`define TANH_LUT_1048 16'h1048
`define TANH_LUT_1050 16'h1050
`define TANH_LUT_1058 16'h1058
`define TANH_LUT_1060 16'h1060
`define TANH_LUT_1068 16'h1068
`define TANH_LUT_1070 16'h1070
`define TANH_LUT_1078 16'h1078
`define TANH_LUT_1080 16'h1080
`define TANH_LUT_1088 16'h1088
`define TANH_LUT_1090 16'h1090
`define TANH_LUT_1098 16'h1098
`define TANH_LUT_10A0 16'h10A0
`define TANH_LUT_10A8 16'h10A8
`define TANH_LUT_10B0 16'h10B0
`define TANH_LUT_10B8 16'h10B8
`define TANH_LUT_10C0 16'h10C0
`define TANH_LUT_10C8 16'h10C8
`define TANH_LUT_10D0 16'h10D0
`define TANH_LUT_10D8 16'h10D8
`define TANH_LUT_10E0 16'h10E0
`define TANH_LUT_10E8 16'h10E8
`define TANH_LUT_10F0 16'h10F0
`define TANH_LUT_10F8 16'h10F8
`define TANH_LUT_1100 16'h1100
`define TANH_LUT_1108 16'h1108
`define TANH_LUT_1110 16'h1110
`define TANH_LUT_1118 16'h1118
`define TANH_LUT_1120 16'h1120
`define TANH_LUT_1128 16'h1128
`define TANH_LUT_1130 16'h1130
`define TANH_LUT_1138 16'h1138
`define TANH_LUT_1140 16'h1140
`define TANH_LUT_1148 16'h1148
`define TANH_LUT_1150 16'h1150
`define TANH_LUT_1158 16'h1158
`define TANH_LUT_1160 16'h1160
`define TANH_LUT_1168 16'h1168
`define TANH_LUT_1170 16'h1170
`define TANH_LUT_1178 16'h1178
`define TANH_LUT_1180 16'h1180
`define TANH_LUT_1188 16'h1188
`define TANH_LUT_1190 16'h1190
`define TANH_LUT_1198 16'h1198
`define TANH_LUT_11A0 16'h11A0
`define TANH_LUT_11A8 16'h11A8
`define TANH_LUT_11B0 16'h11B0
`define TANH_LUT_11B8 16'h11B8
`define TANH_LUT_11C0 16'h11C0
`define TANH_LUT_11C8 16'h11C8
`define TANH_LUT_11D0 16'h11D0
`define TANH_LUT_11D8 16'h11D8
`define TANH_LUT_11E0 16'h11E0
`define TANH_LUT_11E8 16'h11E8
`define TANH_LUT_11F0 16'h11F0
`define TANH_LUT_11F8 16'h11F8
`define TANH_LUT_1200 16'h1200
`define TANH_LUT_1208 16'h1208
`define TANH_LUT_1210 16'h1210
`define TANH_LUT_1218 16'h1218
`define TANH_LUT_1220 16'h1220
`define TANH_LUT_1228 16'h1228
`define TANH_LUT_1230 16'h1230
`define TANH_LUT_1238 16'h1238
`define TANH_LUT_1240 16'h1240
`define TANH_LUT_1248 16'h1248
`define TANH_LUT_1250 16'h1250
`define TANH_LUT_1258 16'h1258
`define TANH_LUT_1260 16'h1260
`define TANH_LUT_1268 16'h1268
`define TANH_LUT_1270 16'h1270
`define TANH_LUT_1278 16'h1278
`define TANH_LUT_1280 16'h1280
`define TANH_LUT_1288 16'h1288
`define TANH_LUT_1290 16'h1290
`define TANH_LUT_1298 16'h1298
`define TANH_LUT_12A0 16'h12A0
`define TANH_LUT_12A8 16'h12A8
`define TANH_LUT_12B0 16'h12B0
`define TANH_LUT_12B8 16'h12B8
`define TANH_LUT_12C0 16'h12C0
`define TANH_LUT_12C8 16'h12C8
`define TANH_LUT_12D0 16'h12D0
`define TANH_LUT_12D8 16'h12D8
`define TANH_LUT_12E0 16'h12E0
`define TANH_LUT_12E8 16'h12E8
`define TANH_LUT_12F0 16'h12F0
`define TANH_LUT_12F8 16'h12F8
`define TANH_LUT_1300 16'h1300
`define TANH_LUT_1308 16'h1308
`define TANH_LUT_1310 16'h1310
`define TANH_LUT_1318 16'h1318
`define TANH_LUT_1320 16'h1320
`define TANH_LUT_1328 16'h1328
`define TANH_LUT_1330 16'h1330
`define TANH_LUT_1338 16'h1338
`define TANH_LUT_1340 16'h1340
`define TANH_LUT_1348 16'h1348
`define TANH_LUT_1350 16'h1350
`define TANH_LUT_1358 16'h1358
`define TANH_LUT_1360 16'h1360
`define TANH_LUT_1368 16'h1368
`define TANH_LUT_1370 16'h1370
`define TANH_LUT_1378 16'h1378
`define TANH_LUT_1380 16'h1380
`define TANH_LUT_1388 16'h1388
`define TANH_LUT_1390 16'h1390
`define TANH_LUT_1398 16'h1398
`define TANH_LUT_13A0 16'h13A0
`define TANH_LUT_13A8 16'h13A8
`define TANH_LUT_13B0 16'h13B0
`define TANH_LUT_13B8 16'h13B8
`define TANH_LUT_13C0 16'h13C0
`define TANH_LUT_13C8 16'h13C8
`define TANH_LUT_13D0 16'h13D0
`define TANH_LUT_13D8 16'h13D8
`define TANH_LUT_13E0 16'h13E0
`define TANH_LUT_13E8 16'h13E8
`define TANH_LUT_13F0 16'h13F0
`define TANH_LUT_13F8 16'h13F8
`define TANH_LUT_1400 16'h1400
`define TANH_LUT_1408 16'h1408
`define TANH_LUT_1410 16'h1410
`define TANH_LUT_1418 16'h1418
`define TANH_LUT_1420 16'h1420
`define TANH_LUT_1428 16'h1428
`define TANH_LUT_1430 16'h1430
`define TANH_LUT_1438 16'h1438
`define TANH_LUT_1440 16'h1440
`define TANH_LUT_1448 16'h1448
`define TANH_LUT_1450 16'h1450
`define TANH_LUT_1458 16'h1458
`define TANH_LUT_1460 16'h1460
`define TANH_LUT_1468 16'h1468
`define TANH_LUT_1470 16'h1470
`define TANH_LUT_1478 16'h1478
`define TANH_LUT_1480 16'h1480
`define TANH_LUT_1488 16'h1488
`define TANH_LUT_1490 16'h1490
`define TANH_LUT_1498 16'h1498
`define TANH_LUT_14A0 16'h14A0
`define TANH_LUT_14A8 16'h14A8
`define TANH_LUT_14B0 16'h14B0
`define TANH_LUT_14B8 16'h14B8
`define TANH_LUT_14C0 16'h14C0
`define TANH_LUT_14C8 16'h14C8
`define TANH_LUT_14D0 16'h14D0
`define TANH_LUT_14D8 16'h14D8
`define TANH_LUT_14E0 16'h14E0
`define TANH_LUT_14E8 16'h14E8
`define TANH_LUT_14F0 16'h14F0
`define TANH_LUT_14F8 16'h14F8
`define TANH_LUT_1500 16'h1500
`define TANH_LUT_1508 16'h1508
`define TANH_LUT_1510 16'h1510
`define TANH_LUT_1518 16'h1518
`define TANH_LUT_1520 16'h1520
`define TANH_LUT_1528 16'h1528
`define TANH_LUT_1530 16'h1530
`define TANH_LUT_1538 16'h1538
`define TANH_LUT_1540 16'h1540
`define TANH_LUT_1548 16'h1548
`define TANH_LUT_1550 16'h1550
`define TANH_LUT_1558 16'h1558
`define TANH_LUT_1560 16'h1560
`define TANH_LUT_1568 16'h1568
`define TANH_LUT_1570 16'h1570
`define TANH_LUT_1578 16'h1578
`define TANH_LUT_1580 16'h1580
`define TANH_LUT_1588 16'h1588
`define TANH_LUT_1590 16'h1590
`define TANH_LUT_1598 16'h1598
`define TANH_LUT_15A0 16'h15A0
`define TANH_LUT_15A8 16'h15A8
`define TANH_LUT_15B0 16'h15B0
`define TANH_LUT_15B8 16'h15B8
`define TANH_LUT_15C0 16'h15C0
`define TANH_LUT_15C8 16'h15C8
`define TANH_LUT_15D0 16'h15D0
`define TANH_LUT_15D8 16'h15D8
`define TANH_LUT_15E0 16'h15E0
`define TANH_LUT_15E8 16'h15E8
`define TANH_LUT_15F0 16'h15F0
`define TANH_LUT_15F8 16'h15F8
`define TANH_LUT_1600 16'h1600
`define TANH_LUT_1608 16'h1608
`define TANH_LUT_1610 16'h1610
`define TANH_LUT_1618 16'h1618
`define TANH_LUT_1620 16'h1620
`define TANH_LUT_1628 16'h1628
`define TANH_LUT_1630 16'h1630
`define TANH_LUT_1638 16'h1638
`define TANH_LUT_1640 16'h1640
`define TANH_LUT_1648 16'h1648
`define TANH_LUT_1650 16'h1650
`define TANH_LUT_1658 16'h1658
`define TANH_LUT_1660 16'h1660
`define TANH_LUT_1668 16'h1668
`define TANH_LUT_1670 16'h1670
`define TANH_LUT_1678 16'h1678
`define TANH_LUT_1680 16'h1680
`define TANH_LUT_1688 16'h1688
`define TANH_LUT_1690 16'h1690
`define TANH_LUT_1698 16'h1698
`define TANH_LUT_16A0 16'h16A0
`define TANH_LUT_16A8 16'h16A8
`define TANH_LUT_16B0 16'h16B0
`define TANH_LUT_16B8 16'h16B8
`define TANH_LUT_16C0 16'h16C0
`define TANH_LUT_16C8 16'h16C8
`define TANH_LUT_16D0 16'h16D0
`define TANH_LUT_16D8 16'h16D8
`define TANH_LUT_16E0 16'h16E0
`define TANH_LUT_16E8 16'h16E8
`define TANH_LUT_16F0 16'h16F0
`define TANH_LUT_16F8 16'h16F8
`define TANH_LUT_1700 16'h1700
`define TANH_LUT_1708 16'h1708
`define TANH_LUT_1710 16'h1710
`define TANH_LUT_1718 16'h1718
`define TANH_LUT_1720 16'h1720
`define TANH_LUT_1728 16'h1728
`define TANH_LUT_1730 16'h1730
`define TANH_LUT_1738 16'h1738
`define TANH_LUT_1740 16'h1740
`define TANH_LUT_1748 16'h1748
`define TANH_LUT_1750 16'h1750
`define TANH_LUT_1758 16'h1758
`define TANH_LUT_1760 16'h1760
`define TANH_LUT_1768 16'h1768
`define TANH_LUT_1770 16'h1770
`define TANH_LUT_1778 16'h1778
`define TANH_LUT_1780 16'h1780
`define TANH_LUT_1788 16'h1788
`define TANH_LUT_1790 16'h1790
`define TANH_LUT_1798 16'h1798
`define TANH_LUT_17A0 16'h17A0
`define TANH_LUT_17A8 16'h17A8
`define TANH_LUT_17B0 16'h17B0
`define TANH_LUT_17B8 16'h17B8
`define TANH_LUT_17C0 16'h17C0
`define TANH_LUT_17C8 16'h17C8
`define TANH_LUT_17D0 16'h17D0
`define TANH_LUT_17D8 16'h17D8
`define TANH_LUT_17E0 16'h17E0
`define TANH_LUT_17E8 16'h17E8
`define TANH_LUT_17F0 16'h17F0
`define TANH_LUT_17F8 16'h17F8
`define TANH_LUT_1800 16'h1800
`define TANH_LUT_1808 16'h1808
`define TANH_LUT_1810 16'h1810
`define TANH_LUT_1818 16'h1818
`define TANH_LUT_1820 16'h1820
`define TANH_LUT_1828 16'h1828
`define TANH_LUT_1830 16'h1830
`define TANH_LUT_1838 16'h1838
`define TANH_LUT_1840 16'h1840
`define TANH_LUT_1848 16'h1848
`define TANH_LUT_1850 16'h1850
`define TANH_LUT_1858 16'h1858
`define TANH_LUT_1860 16'h1860
`define TANH_LUT_1868 16'h1868
`define TANH_LUT_1870 16'h1870
`define TANH_LUT_1878 16'h1878
`define TANH_LUT_1880 16'h1880
`define TANH_LUT_1888 16'h1888
`define TANH_LUT_1890 16'h1890
`define TANH_LUT_1898 16'h1898
`define TANH_LUT_18A0 16'h18A0
`define TANH_LUT_18A8 16'h18A8
`define TANH_LUT_18B0 16'h18B0
`define TANH_LUT_18B8 16'h18B8
`define TANH_LUT_18C0 16'h18C0
`define TANH_LUT_18C8 16'h18C8
`define TANH_LUT_18D0 16'h18D0
`define TANH_LUT_18D8 16'h18D8
`define TANH_LUT_18E0 16'h18E0
`define TANH_LUT_18E8 16'h18E8
`define TANH_LUT_18F0 16'h18F0
`define TANH_LUT_18F8 16'h18F8
`define TANH_LUT_1900 16'h1900
`define TANH_LUT_1908 16'h1908
`define TANH_LUT_1910 16'h1910
`define TANH_LUT_1918 16'h1918
`define TANH_LUT_1920 16'h1920
`define TANH_LUT_1928 16'h1928
`define TANH_LUT_1930 16'h1930
`define TANH_LUT_1938 16'h1938
`define TANH_LUT_1940 16'h1940
`define TANH_LUT_1948 16'h1948
`define TANH_LUT_1950 16'h1950
`define TANH_LUT_1958 16'h1958
`define TANH_LUT_1960 16'h1960
`define TANH_LUT_1968 16'h1968
`define TANH_LUT_1970 16'h1970
`define TANH_LUT_1978 16'h1978
`define TANH_LUT_1980 16'h1980
`define TANH_LUT_1988 16'h1988
`define TANH_LUT_1990 16'h1990
`define TANH_LUT_1998 16'h1998
`define TANH_LUT_19A0 16'h19A0
`define TANH_LUT_19A8 16'h19A8
`define TANH_LUT_19B0 16'h19B0
`define TANH_LUT_19B8 16'h19B8
`define TANH_LUT_19C0 16'h19C0
`define TANH_LUT_19C8 16'h19C8
`define TANH_LUT_19D0 16'h19D0
`define TANH_LUT_19D8 16'h19D8
`define TANH_LUT_19E0 16'h19E0
`define TANH_LUT_19E8 16'h19E8
`define TANH_LUT_19F0 16'h19F0
`define TANH_LUT_19F8 16'h19F8
`define TANH_LUT_1A00 16'h1A00
`define TANH_LUT_1A08 16'h1A08
`define TANH_LUT_1A10 16'h1A10
`define TANH_LUT_1A18 16'h1A18
`define TANH_LUT_1A20 16'h1A20
`define TANH_LUT_1A28 16'h1A28
`define TANH_LUT_1A30 16'h1A30
`define TANH_LUT_1A38 16'h1A38
`define TANH_LUT_1A40 16'h1A40
`define TANH_LUT_1A48 16'h1A48
`define TANH_LUT_1A50 16'h1A50
`define TANH_LUT_1A58 16'h1A58
`define TANH_LUT_1A60 16'h1A60
`define TANH_LUT_1A68 16'h1A68
`define TANH_LUT_1A70 16'h1A70
`define TANH_LUT_1A78 16'h1A78
`define TANH_LUT_1A80 16'h1A80
`define TANH_LUT_1A88 16'h1A88
`define TANH_LUT_1A90 16'h1A90
`define TANH_LUT_1A98 16'h1A98
`define TANH_LUT_1AA0 16'h1AA0
`define TANH_LUT_1AA8 16'h1AA8
`define TANH_LUT_1AB0 16'h1AB0
`define TANH_LUT_1AB8 16'h1AB8
`define TANH_LUT_1AC0 16'h1AC0
`define TANH_LUT_1AC8 16'h1AC8
`define TANH_LUT_1AD0 16'h1AD0
`define TANH_LUT_1AD8 16'h1AD8
`define TANH_LUT_1AE0 16'h1AE0
`define TANH_LUT_1AE8 16'h1AE8
`define TANH_LUT_1AF0 16'h1AF0
`define TANH_LUT_1AF8 16'h1AF8
`define TANH_LUT_1B00 16'h1B00
`define TANH_LUT_1B08 16'h1B08
`define TANH_LUT_1B10 16'h1B10
`define TANH_LUT_1B18 16'h1B18
`define TANH_LUT_1B20 16'h1B20
`define TANH_LUT_1B28 16'h1B28
`define TANH_LUT_1B30 16'h1B30
`define TANH_LUT_1B38 16'h1B38
`define TANH_LUT_1B40 16'h1B40
`define TANH_LUT_1B48 16'h1B48
`define TANH_LUT_1B50 16'h1B50
`define TANH_LUT_1B58 16'h1B58
`define TANH_LUT_1B60 16'h1B60
`define TANH_LUT_1B68 16'h1B68
`define TANH_LUT_1B70 16'h1B70
`define TANH_LUT_1B78 16'h1B78
`define TANH_LUT_1B80 16'h1B80
`define TANH_LUT_1B88 16'h1B88
`define TANH_LUT_1B90 16'h1B90
`define TANH_LUT_1B98 16'h1B98
`define TANH_LUT_1BA0 16'h1BA0
`define TANH_LUT_1BA8 16'h1BA8
`define TANH_LUT_1BB0 16'h1BB0
`define TANH_LUT_1BB8 16'h1BB8
`define TANH_LUT_1BC0 16'h1BC0
`define TANH_LUT_1BC8 16'h1BC8
`define TANH_LUT_1BD0 16'h1BD0
`define TANH_LUT_1BD8 16'h1BD8
`define TANH_LUT_1BE0 16'h1BE0
`define TANH_LUT_1BE8 16'h1BE8
`define TANH_LUT_1BF0 16'h1BF0
`define TANH_LUT_1BF8 16'h1BF8
`define TANH_LUT_1C00 16'h1C00
`define TANH_LUT_1C08 16'h1C08
`define TANH_LUT_1C10 16'h1C10
`define TANH_LUT_1C18 16'h1C18
`define TANH_LUT_1C20 16'h1C20
`define TANH_LUT_1C28 16'h1C28
`define TANH_LUT_1C30 16'h1C30
`define TANH_LUT_1C38 16'h1C38
`define TANH_LUT_1C40 16'h1C40
`define TANH_LUT_1C48 16'h1C48
`define TANH_LUT_1C50 16'h1C50
`define TANH_LUT_1C58 16'h1C58
`define TANH_LUT_1C60 16'h1C60
`define TANH_LUT_1C68 16'h1C68
`define TANH_LUT_1C70 16'h1C70
`define TANH_LUT_1C78 16'h1C78
`define TANH_LUT_1C80 16'h1C80
`define TANH_LUT_1C88 16'h1C88
`define TANH_LUT_1C90 16'h1C90
`define TANH_LUT_1C98 16'h1C98
`define TANH_LUT_1CA0 16'h1CA0
`define TANH_LUT_1CA8 16'h1CA8
`define TANH_LUT_1CB0 16'h1CB0
`define TANH_LUT_1CB8 16'h1CB8
`define TANH_LUT_1CC0 16'h1CC0
`define TANH_LUT_1CC8 16'h1CC8
`define TANH_LUT_1CD0 16'h1CD0
`define TANH_LUT_1CD8 16'h1CD8
`define TANH_LUT_1CE0 16'h1CE0
`define TANH_LUT_1CE8 16'h1CE8
`define TANH_LUT_1CF0 16'h1CF0
`define TANH_LUT_1CF8 16'h1CF8
`define TANH_LUT_1D00 16'h1D00
`define TANH_LUT_1D08 16'h1D08
`define TANH_LUT_1D10 16'h1D10
`define TANH_LUT_1D18 16'h1D18
`define TANH_LUT_1D20 16'h1D20
`define TANH_LUT_1D28 16'h1D28
`define TANH_LUT_1D30 16'h1D30
`define TANH_LUT_1D38 16'h1D38
`define TANH_LUT_1D40 16'h1D40
`define TANH_LUT_1D48 16'h1D48
`define TANH_LUT_1D50 16'h1D50
`define TANH_LUT_1D58 16'h1D58
`define TANH_LUT_1D60 16'h1D60
`define TANH_LUT_1D68 16'h1D68
`define TANH_LUT_1D70 16'h1D70
`define TANH_LUT_1D78 16'h1D78
`define TANH_LUT_1D80 16'h1D80
`define TANH_LUT_1D88 16'h1D88
`define TANH_LUT_1D90 16'h1D90
`define TANH_LUT_1D98 16'h1D98
`define TANH_LUT_1DA0 16'h1DA0
`define TANH_LUT_1DA8 16'h1DA8
`define TANH_LUT_1DB0 16'h1DB0
`define TANH_LUT_1DB8 16'h1DB8
`define TANH_LUT_1DC0 16'h1DC0
`define TANH_LUT_1DC8 16'h1DC8
`define TANH_LUT_1DD0 16'h1DD0
`define TANH_LUT_1DD8 16'h1DD8
`define TANH_LUT_1DE0 16'h1DE0
`define TANH_LUT_1DE8 16'h1DE8
`define TANH_LUT_1DF0 16'h1DF0
`define TANH_LUT_1DF8 16'h1DF8
`define TANH_LUT_1E00 16'h1E00
`define TANH_LUT_1E08 16'h1E08
`define TANH_LUT_1E10 16'h1E10
`define TANH_LUT_1E18 16'h1E18
`define TANH_LUT_1E20 16'h1E20
`define TANH_LUT_1E28 16'h1E28
`define TANH_LUT_1E30 16'h1E30
`define TANH_LUT_1E38 16'h1E38
`define TANH_LUT_1E40 16'h1E40
`define TANH_LUT_1E48 16'h1E48
`define TANH_LUT_1E50 16'h1E50
`define TANH_LUT_1E58 16'h1E58
`define TANH_LUT_1E60 16'h1E60
`define TANH_LUT_1E68 16'h1E68
`define TANH_LUT_1E70 16'h1E70
`define TANH_LUT_1E78 16'h1E78
`define TANH_LUT_1E80 16'h1E80
`define TANH_LUT_1E88 16'h1E88
`define TANH_LUT_1E90 16'h1E90
`define TANH_LUT_1E98 16'h1E98
`define TANH_LUT_1EA0 16'h1EA0
`define TANH_LUT_1EA8 16'h1EA8
`define TANH_LUT_1EB0 16'h1EB0
`define TANH_LUT_1EB8 16'h1EB8
`define TANH_LUT_1EC0 16'h1EC0
`define TANH_LUT_1EC8 16'h1EC8
`define TANH_LUT_1ED0 16'h1ED0
`define TANH_LUT_1ED8 16'h1ED8
`define TANH_LUT_1EE0 16'h1EE0
`define TANH_LUT_1EE8 16'h1EE8
`define TANH_LUT_1EF0 16'h1EF0
`define TANH_LUT_1EF8 16'h1EF8
`define TANH_LUT_1F00 16'h1F00
`define TANH_LUT_1F08 16'h1F08
`define TANH_LUT_1F10 16'h1F10
`define TANH_LUT_1F18 16'h1F18
`define TANH_LUT_1F20 16'h1F20
`define TANH_LUT_1F28 16'h1F28
`define TANH_LUT_1F30 16'h1F30
`define TANH_LUT_1F38 16'h1F38
`define TANH_LUT_1F40 16'h1F40
`define TANH_LUT_1F48 16'h1F48
`define TANH_LUT_1F50 16'h1F50
`define TANH_LUT_1F58 16'h1F58
`define TANH_LUT_1F60 16'h1F60
`define TANH_LUT_1F68 16'h1F68
`define TANH_LUT_1F70 16'h1F70
`define TANH_LUT_1F78 16'h1F78
`define TANH_LUT_1F80 16'h1F80
`define TANH_LUT_1F88 16'h1F88
`define TANH_LUT_1F90 16'h1F90
`define TANH_LUT_1F98 16'h1F98
`define TANH_LUT_1FA0 16'h1FA0
`define TANH_LUT_1FA8 16'h1FA8
`define TANH_LUT_1FB0 16'h1FB0
`define TANH_LUT_1FB8 16'h1FB8
`define TANH_LUT_1FC0 16'h1FC0
`define TANH_LUT_1FC8 16'h1FC8
`define TANH_LUT_1FD0 16'h1FD0
`define TANH_LUT_1FD8 16'h1FD8
`define TANH_LUT_1FE0 16'h1FE0
`define TANH_LUT_1FE8 16'h1FE8
`define TANH_LUT_1FF0 16'h1FF0
`define TANH_LUT_1FF8 16'h1FF8
`define TANH_LUT_2000 16'h2000
`define TANH_LUT_2008 16'h2008
`define TANH_LUT_2010 16'h2010
`define TANH_LUT_2018 16'h2018
`define TANH_LUT_2020 16'h2020
`define TANH_LUT_2028 16'h2028
`define TANH_LUT_2030 16'h2030
`define TANH_LUT_2038 16'h2038
`define TANH_LUT_2040 16'h2040
`define TANH_LUT_2048 16'h2048
`define TANH_LUT_2050 16'h2050
`define TANH_LUT_2058 16'h2058
`define TANH_LUT_2060 16'h2060
`define TANH_LUT_2068 16'h2068
`define TANH_LUT_2070 16'h2070
`define TANH_LUT_2078 16'h2078
`define TANH_LUT_2080 16'h2080
`define TANH_LUT_2088 16'h2088
`define TANH_LUT_2090 16'h2090
`define TANH_LUT_2098 16'h2098
`define TANH_LUT_20A0 16'h20A0
`define TANH_LUT_20A8 16'h20A8
`define TANH_LUT_20B0 16'h20B0
`define TANH_LUT_20B8 16'h20B8
`define TANH_LUT_20C0 16'h20C0
`define TANH_LUT_20C8 16'h20C8
`define TANH_LUT_20D0 16'h20D0
`define TANH_LUT_20D8 16'h20D8
`define TANH_LUT_20E0 16'h20E0
`define TANH_LUT_20E8 16'h20E8
`define TANH_LUT_20F0 16'h20F0
`define TANH_LUT_20F8 16'h20F8
`define TANH_LUT_2100 16'h2100
`define TANH_LUT_2108 16'h2108
`define TANH_LUT_2110 16'h2110
`define TANH_LUT_2118 16'h2118
`define TANH_LUT_2120 16'h2120
`define TANH_LUT_2128 16'h2128
`define TANH_LUT_2130 16'h2130
`define TANH_LUT_2138 16'h2138
`define TANH_LUT_2140 16'h2140
`define TANH_LUT_2148 16'h2148
`define TANH_LUT_2150 16'h2150
`define TANH_LUT_2158 16'h2158
`define TANH_LUT_2160 16'h2160
`define TANH_LUT_2168 16'h2168
`define TANH_LUT_2170 16'h2170
`define TANH_LUT_2178 16'h2178
`define TANH_LUT_2180 16'h2180
`define TANH_LUT_2188 16'h2188
`define TANH_LUT_2190 16'h2190
`define TANH_LUT_2198 16'h2198
`define TANH_LUT_21A0 16'h21A0
`define TANH_LUT_21A8 16'h21A8
`define TANH_LUT_21B0 16'h21B0
`define TANH_LUT_21B8 16'h21B8
`define TANH_LUT_21C0 16'h21C0
`define TANH_LUT_21C8 16'h21C8
`define TANH_LUT_21D0 16'h21D0
`define TANH_LUT_21D8 16'h21D8
`define TANH_LUT_21E0 16'h21E0
`define TANH_LUT_21E8 16'h21E8
`define TANH_LUT_21F0 16'h21F0
`define TANH_LUT_21F8 16'h21F8
`define TANH_LUT_2200 16'h2200
`define TANH_LUT_2208 16'h2208
`define TANH_LUT_2210 16'h2210
`define TANH_LUT_2218 16'h2218
`define TANH_LUT_2220 16'h2220
`define TANH_LUT_2228 16'h2228
`define TANH_LUT_2230 16'h2230
`define TANH_LUT_2238 16'h2238
`define TANH_LUT_2240 16'h2240
`define TANH_LUT_2248 16'h2248
`define TANH_LUT_2250 16'h2250
`define TANH_LUT_2258 16'h2258
`define TANH_LUT_2260 16'h2260
`define TANH_LUT_2268 16'h2268
`define TANH_LUT_2270 16'h2270
`define TANH_LUT_2278 16'h2278
`define TANH_LUT_2280 16'h2280
`define TANH_LUT_2288 16'h2288
`define TANH_LUT_2290 16'h2290
`define TANH_LUT_2298 16'h2298
`define TANH_LUT_22A0 16'h22A0
`define TANH_LUT_22A8 16'h22A8
`define TANH_LUT_22B0 16'h22B0
`define TANH_LUT_22B8 16'h22B8
`define TANH_LUT_22C0 16'h22C0
`define TANH_LUT_22C8 16'h22C8
`define TANH_LUT_22D0 16'h22D0
`define TANH_LUT_22D8 16'h22D8
`define TANH_LUT_22E0 16'h22E0
`define TANH_LUT_22E8 16'h22E8
`define TANH_LUT_22F0 16'h22F0
`define TANH_LUT_22F8 16'h22F8
`define TANH_LUT_2300 16'h2300
`define TANH_LUT_2308 16'h2308
`define TANH_LUT_2310 16'h2310
`define TANH_LUT_2318 16'h2318
`define TANH_LUT_2320 16'h2320
`define TANH_LUT_2328 16'h2328
`define TANH_LUT_2330 16'h2330
`define TANH_LUT_2338 16'h2338
`define TANH_LUT_2340 16'h2340
`define TANH_LUT_2348 16'h2348
`define TANH_LUT_2350 16'h2350
`define TANH_LUT_2358 16'h2358
`define TANH_LUT_2360 16'h2360
`define TANH_LUT_2368 16'h2368
`define TANH_LUT_2370 16'h2370
`define TANH_LUT_2378 16'h2378
`define TANH_LUT_2380 16'h2380
`define TANH_LUT_2388 16'h2388
`define TANH_LUT_2390 16'h2390
`define TANH_LUT_2398 16'h2398
`define TANH_LUT_23A0 16'h23A0
`define TANH_LUT_23A8 16'h23A8
`define TANH_LUT_23B0 16'h23B0
`define TANH_LUT_23B8 16'h23B8
`define TANH_LUT_23C0 16'h23C0
`define TANH_LUT_23C8 16'h23C8
`define TANH_LUT_23D0 16'h23D0
`define TANH_LUT_23D8 16'h23D8
`define TANH_LUT_23E0 16'h23E0
`define TANH_LUT_23E8 16'h23E8
`define TANH_LUT_23F0 16'h23F0
`define TANH_LUT_23F8 16'h23F8
`define TANH_LUT_2400 16'h2400
`define TANH_LUT_2408 16'h2408
`define TANH_LUT_2410 16'h2410
`define TANH_LUT_2418 16'h2418
`define TANH_LUT_2420 16'h2420
`define TANH_LUT_2428 16'h2428
`define TANH_LUT_2430 16'h2430
`define TANH_LUT_2438 16'h2438
`define TANH_LUT_2440 16'h2440
`define TANH_LUT_2448 16'h2448
`define TANH_LUT_2450 16'h2450
`define TANH_LUT_2458 16'h2458
`define TANH_LUT_2460 16'h2460
`define TANH_LUT_2468 16'h2468
`define TANH_LUT_2470 16'h2470
`define TANH_LUT_2478 16'h2478
`define TANH_LUT_2480 16'h2480
`define TANH_LUT_2488 16'h2488
`define TANH_LUT_2490 16'h2490
`define TANH_LUT_2498 16'h2498
`define TANH_LUT_24A0 16'h24A0
`define TANH_LUT_24A8 16'h24A8
`define TANH_LUT_24B0 16'h24B0
`define TANH_LUT_24B8 16'h24B8
`define TANH_LUT_24C0 16'h24C0
`define TANH_LUT_24C8 16'h24C8
`define TANH_LUT_24D0 16'h24D0
`define TANH_LUT_24D8 16'h24D8
`define TANH_LUT_24E0 16'h24E0
`define TANH_LUT_24E8 16'h24E8
`define TANH_LUT_24F0 16'h24F0
`define TANH_LUT_24F8 16'h24F8
`define TANH_LUT_2500 16'h2500
`define TANH_LUT_2508 16'h2508
`define TANH_LUT_2510 16'h2510
`define TANH_LUT_2518 16'h2518
`define TANH_LUT_2520 16'h2520
`define TANH_LUT_2528 16'h2528
`define TANH_LUT_2530 16'h2530
`define TANH_LUT_2538 16'h2538
`define TANH_LUT_2540 16'h2540
`define TANH_LUT_2548 16'h2548
`define TANH_LUT_2550 16'h2550
`define TANH_LUT_2558 16'h2558
`define TANH_LUT_2560 16'h2560
`define TANH_LUT_2568 16'h2568
`define TANH_LUT_2570 16'h2570
`define TANH_LUT_2578 16'h2578
`define TANH_LUT_2580 16'h2580
`define TANH_LUT_2588 16'h2588
`define TANH_LUT_2590 16'h2590
`define TANH_LUT_2598 16'h2598
`define TANH_LUT_25A0 16'h25A0
`define TANH_LUT_25A8 16'h25A8
`define TANH_LUT_25B0 16'h25B0
`define TANH_LUT_25B8 16'h25B8
`define TANH_LUT_25C0 16'h25C0
`define TANH_LUT_25C8 16'h25C8
`define TANH_LUT_25D0 16'h25D0
`define TANH_LUT_25D8 16'h25D8
`define TANH_LUT_25E0 16'h25E0
`define TANH_LUT_25E8 16'h25E8
`define TANH_LUT_25F0 16'h25F0
`define TANH_LUT_25F8 16'h25F8
`define TANH_LUT_2600 16'h2600
`define TANH_LUT_2608 16'h2608
`define TANH_LUT_2610 16'h2610
`define TANH_LUT_2618 16'h2618
`define TANH_LUT_2620 16'h2620
`define TANH_LUT_2628 16'h2628
`define TANH_LUT_2630 16'h2630
`define TANH_LUT_2638 16'h2638
`define TANH_LUT_2640 16'h2640
`define TANH_LUT_2648 16'h2648
`define TANH_LUT_2650 16'h2650
`define TANH_LUT_2658 16'h2658
`define TANH_LUT_2660 16'h2660
`define TANH_LUT_2668 16'h2668
`define TANH_LUT_2670 16'h2670
`define TANH_LUT_2678 16'h2678
`define TANH_LUT_2680 16'h2680
`define TANH_LUT_2688 16'h2688
`define TANH_LUT_2690 16'h2690
`define TANH_LUT_2698 16'h2698
`define TANH_LUT_26A0 16'h26A0
`define TANH_LUT_26A8 16'h26A8
`define TANH_LUT_26B0 16'h26B0
`define TANH_LUT_26B8 16'h26B8
`define TANH_LUT_26C0 16'h26C0
`define TANH_LUT_26C8 16'h26C8
`define TANH_LUT_26D0 16'h26D0
`define TANH_LUT_26D8 16'h26D8
`define TANH_LUT_26E0 16'h26E0
`define TANH_LUT_26E8 16'h26E8
`define TANH_LUT_26F0 16'h26F0
`define TANH_LUT_26F8 16'h26F8
`define TANH_LUT_2700 16'h2700
`define TANH_LUT_2708 16'h2708
`define TANH_LUT_2710 16'h2710
`define TANH_LUT_2718 16'h2718
`define TANH_LUT_2720 16'h2720
`define TANH_LUT_2728 16'h2728
`define TANH_LUT_2730 16'h2730
`define TANH_LUT_2738 16'h2738
`define TANH_LUT_2740 16'h2740
`define TANH_LUT_2748 16'h2747
`define TANH_LUT_2750 16'h274F
`define TANH_LUT_2758 16'h2757
`define TANH_LUT_2760 16'h275F
`define TANH_LUT_2768 16'h2767
`define TANH_LUT_2770 16'h276F
`define TANH_LUT_2778 16'h2777
`define TANH_LUT_2780 16'h277F
`define TANH_LUT_2788 16'h2787
`define TANH_LUT_2790 16'h278F
`define TANH_LUT_2798 16'h2797
`define TANH_LUT_27A0 16'h279F
`define TANH_LUT_27A8 16'h27A7
`define TANH_LUT_27B0 16'h27AF
`define TANH_LUT_27B8 16'h27B7
`define TANH_LUT_27C0 16'h27BF
`define TANH_LUT_27C8 16'h27C7
`define TANH_LUT_27D0 16'h27CF
`define TANH_LUT_27D8 16'h27D7
`define TANH_LUT_27E0 16'h27DF
`define TANH_LUT_27E8 16'h27E7
`define TANH_LUT_27F0 16'h27EF
`define TANH_LUT_27F8 16'h27F7
`define TANH_LUT_2800 16'h27FF
`define TANH_LUT_2808 16'h2808
`define TANH_LUT_2810 16'h2810
`define TANH_LUT_2818 16'h2818
`define TANH_LUT_2820 16'h2820
`define TANH_LUT_2828 16'h2828
`define TANH_LUT_2830 16'h2830
`define TANH_LUT_2838 16'h2838
`define TANH_LUT_2840 16'h2840
`define TANH_LUT_2848 16'h2848
`define TANH_LUT_2850 16'h2850
`define TANH_LUT_2858 16'h2858
`define TANH_LUT_2860 16'h2860
`define TANH_LUT_2868 16'h2868
`define TANH_LUT_2870 16'h2870
`define TANH_LUT_2878 16'h2878
`define TANH_LUT_2880 16'h2880
`define TANH_LUT_2888 16'h2888
`define TANH_LUT_2890 16'h2890
`define TANH_LUT_2898 16'h2897
`define TANH_LUT_28A0 16'h289F
`define TANH_LUT_28A8 16'h28A7
`define TANH_LUT_28B0 16'h28AF
`define TANH_LUT_28B8 16'h28B7
`define TANH_LUT_28C0 16'h28BF
`define TANH_LUT_28C8 16'h28C7
`define TANH_LUT_28D0 16'h28CF
`define TANH_LUT_28D8 16'h28D7
`define TANH_LUT_28E0 16'h28DF
`define TANH_LUT_28E8 16'h28E7
`define TANH_LUT_28F0 16'h28EF
`define TANH_LUT_28F8 16'h28F7
`define TANH_LUT_2900 16'h28FF
`define TANH_LUT_2908 16'h2907
`define TANH_LUT_2910 16'h290F
`define TANH_LUT_2918 16'h2917
`define TANH_LUT_2920 16'h291F
`define TANH_LUT_2928 16'h2927
`define TANH_LUT_2930 16'h292F
`define TANH_LUT_2938 16'h2937
`define TANH_LUT_2940 16'h293F
`define TANH_LUT_2948 16'h2947
`define TANH_LUT_2950 16'h294F
`define TANH_LUT_2958 16'h2957
`define TANH_LUT_2960 16'h295F
`define TANH_LUT_2968 16'h2967
`define TANH_LUT_2970 16'h296F
`define TANH_LUT_2978 16'h2977
`define TANH_LUT_2980 16'h297F
`define TANH_LUT_2988 16'h2987
`define TANH_LUT_2990 16'h298F
`define TANH_LUT_2998 16'h2997
`define TANH_LUT_29A0 16'h299F
`define TANH_LUT_29A8 16'h29A7
`define TANH_LUT_29B0 16'h29AF
`define TANH_LUT_29B8 16'h29B7
`define TANH_LUT_29C0 16'h29BF
`define TANH_LUT_29C8 16'h29C7
`define TANH_LUT_29D0 16'h29CF
`define TANH_LUT_29D8 16'h29D7
`define TANH_LUT_29E0 16'h29DF
`define TANH_LUT_29E8 16'h29E7
`define TANH_LUT_29F0 16'h29EF
`define TANH_LUT_29F8 16'h29F7
`define TANH_LUT_2A00 16'h29FF
`define TANH_LUT_2A08 16'h2A07
`define TANH_LUT_2A10 16'h2A0F
`define TANH_LUT_2A18 16'h2A17
`define TANH_LUT_2A20 16'h2A1F
`define TANH_LUT_2A28 16'h2A27
`define TANH_LUT_2A30 16'h2A2F
`define TANH_LUT_2A38 16'h2A37
`define TANH_LUT_2A40 16'h2A3F
`define TANH_LUT_2A48 16'h2A47
`define TANH_LUT_2A50 16'h2A4F
`define TANH_LUT_2A58 16'h2A57
`define TANH_LUT_2A60 16'h2A5F
`define TANH_LUT_2A68 16'h2A67
`define TANH_LUT_2A70 16'h2A6F
`define TANH_LUT_2A78 16'h2A77
`define TANH_LUT_2A80 16'h2A7F
`define TANH_LUT_2A88 16'h2A87
`define TANH_LUT_2A90 16'h2A8F
`define TANH_LUT_2A98 16'h2A97
`define TANH_LUT_2AA0 16'h2A9E
`define TANH_LUT_2AA8 16'h2AA6
`define TANH_LUT_2AB0 16'h2AAE
`define TANH_LUT_2AB8 16'h2AB6
`define TANH_LUT_2AC0 16'h2ABE
`define TANH_LUT_2AC8 16'h2AC6
`define TANH_LUT_2AD0 16'h2ACE
`define TANH_LUT_2AD8 16'h2AD6
`define TANH_LUT_2AE0 16'h2ADE
`define TANH_LUT_2AE8 16'h2AE6
`define TANH_LUT_2AF0 16'h2AEE
`define TANH_LUT_2AF8 16'h2AF6
`define TANH_LUT_2B00 16'h2AFE
`define TANH_LUT_2B08 16'h2B06
`define TANH_LUT_2B10 16'h2B0E
`define TANH_LUT_2B18 16'h2B16
`define TANH_LUT_2B20 16'h2B1E
`define TANH_LUT_2B28 16'h2B26
`define TANH_LUT_2B30 16'h2B2E
`define TANH_LUT_2B38 16'h2B36
`define TANH_LUT_2B40 16'h2B3E
`define TANH_LUT_2B48 16'h2B46
`define TANH_LUT_2B50 16'h2B4E
`define TANH_LUT_2B58 16'h2B56
`define TANH_LUT_2B60 16'h2B5E
`define TANH_LUT_2B68 16'h2B66
`define TANH_LUT_2B70 16'h2B6E
`define TANH_LUT_2B78 16'h2B76
`define TANH_LUT_2B80 16'h2B7E
`define TANH_LUT_2B88 16'h2B86
`define TANH_LUT_2B90 16'h2B8E
`define TANH_LUT_2B98 16'h2B96
`define TANH_LUT_2BA0 16'h2B9E
`define TANH_LUT_2BA8 16'h2BA6
`define TANH_LUT_2BB0 16'h2BAE
`define TANH_LUT_2BB8 16'h2BB6
`define TANH_LUT_2BC0 16'h2BBE
`define TANH_LUT_2BC8 16'h2BC6
`define TANH_LUT_2BD0 16'h2BCE
`define TANH_LUT_2BD8 16'h2BD5
`define TANH_LUT_2BE0 16'h2BDD
`define TANH_LUT_2BE8 16'h2BE5
`define TANH_LUT_2BF0 16'h2BED
`define TANH_LUT_2BF8 16'h2BF5
`define TANH_LUT_2C00 16'h2BFD
`define TANH_LUT_2C08 16'h2C07
`define TANH_LUT_2C10 16'h2C0F
`define TANH_LUT_2C18 16'h2C17
`define TANH_LUT_2C20 16'h2C1F
`define TANH_LUT_2C28 16'h2C27
`define TANH_LUT_2C30 16'h2C2E
`define TANH_LUT_2C38 16'h2C36
`define TANH_LUT_2C40 16'h2C3E
`define TANH_LUT_2C48 16'h2C46
`define TANH_LUT_2C50 16'h2C4E
`define TANH_LUT_2C58 16'h2C56
`define TANH_LUT_2C60 16'h2C5E
`define TANH_LUT_2C68 16'h2C66
`define TANH_LUT_2C70 16'h2C6E
`define TANH_LUT_2C78 16'h2C76
`define TANH_LUT_2C80 16'h2C7E
`define TANH_LUT_2C88 16'h2C86
`define TANH_LUT_2C90 16'h2C8E
`define TANH_LUT_2C98 16'h2C96
`define TANH_LUT_2CA0 16'h2C9E
`define TANH_LUT_2CA8 16'h2CA6
`define TANH_LUT_2CB0 16'h2CAE
`define TANH_LUT_2CB8 16'h2CB6
`define TANH_LUT_2CC0 16'h2CBE
`define TANH_LUT_2CC8 16'h2CC6
`define TANH_LUT_2CD0 16'h2CCE
`define TANH_LUT_2CD8 16'h2CD6
`define TANH_LUT_2CE0 16'h2CDE
`define TANH_LUT_2CE8 16'h2CE6
`define TANH_LUT_2CF0 16'h2CED
`define TANH_LUT_2CF8 16'h2CF5
`define TANH_LUT_2D00 16'h2CFD
`define TANH_LUT_2D08 16'h2D05
`define TANH_LUT_2D10 16'h2D0D
`define TANH_LUT_2D18 16'h2D15
`define TANH_LUT_2D20 16'h2D1D
`define TANH_LUT_2D28 16'h2D25
`define TANH_LUT_2D30 16'h2D2D
`define TANH_LUT_2D38 16'h2D35
`define TANH_LUT_2D40 16'h2D3D
`define TANH_LUT_2D48 16'h2D45
`define TANH_LUT_2D50 16'h2D4D
`define TANH_LUT_2D58 16'h2D55
`define TANH_LUT_2D60 16'h2D5D
`define TANH_LUT_2D68 16'h2D65
`define TANH_LUT_2D70 16'h2D6D
`define TANH_LUT_2D78 16'h2D75
`define TANH_LUT_2D80 16'h2D7D
`define TANH_LUT_2D88 16'h2D84
`define TANH_LUT_2D90 16'h2D8C
`define TANH_LUT_2D98 16'h2D94
`define TANH_LUT_2DA0 16'h2D9C
`define TANH_LUT_2DA8 16'h2DA4
`define TANH_LUT_2DB0 16'h2DAC
`define TANH_LUT_2DB8 16'h2DB4
`define TANH_LUT_2DC0 16'h2DBC
`define TANH_LUT_2DC8 16'h2DC4
`define TANH_LUT_2DD0 16'h2DCC
`define TANH_LUT_2DD8 16'h2DD4
`define TANH_LUT_2DE0 16'h2DDC
`define TANH_LUT_2DE8 16'h2DE4
`define TANH_LUT_2DF0 16'h2DEC
`define TANH_LUT_2DF8 16'h2DF4
`define TANH_LUT_2E00 16'h2DFC
`define TANH_LUT_2E08 16'h2E03
`define TANH_LUT_2E10 16'h2E0B
`define TANH_LUT_2E18 16'h2E13
`define TANH_LUT_2E20 16'h2E1B
`define TANH_LUT_2E28 16'h2E23
`define TANH_LUT_2E30 16'h2E2B
`define TANH_LUT_2E38 16'h2E33
`define TANH_LUT_2E40 16'h2E3B
`define TANH_LUT_2E48 16'h2E43
`define TANH_LUT_2E50 16'h2E4B
`define TANH_LUT_2E58 16'h2E53
`define TANH_LUT_2E60 16'h2E5B
`define TANH_LUT_2E68 16'h2E63
`define TANH_LUT_2E70 16'h2E6A
`define TANH_LUT_2E78 16'h2E72
`define TANH_LUT_2E80 16'h2E7A
`define TANH_LUT_2E88 16'h2E82
`define TANH_LUT_2E90 16'h2E8A
`define TANH_LUT_2E98 16'h2E92
`define TANH_LUT_2EA0 16'h2E9A
`define TANH_LUT_2EA8 16'h2EA2
`define TANH_LUT_2EB0 16'h2EAA
`define TANH_LUT_2EB8 16'h2EB2
`define TANH_LUT_2EC0 16'h2EBA
`define TANH_LUT_2EC8 16'h2EC2
`define TANH_LUT_2ED0 16'h2EC9
`define TANH_LUT_2ED8 16'h2ED1
`define TANH_LUT_2EE0 16'h2ED9
`define TANH_LUT_2EE8 16'h2EE1
`define TANH_LUT_2EF0 16'h2EE9
`define TANH_LUT_2EF8 16'h2EF1
`define TANH_LUT_2F00 16'h2EF9
`define TANH_LUT_2F08 16'h2F01
`define TANH_LUT_2F10 16'h2F09
`define TANH_LUT_2F18 16'h2F11
`define TANH_LUT_2F20 16'h2F19
`define TANH_LUT_2F28 16'h2F20
`define TANH_LUT_2F30 16'h2F28
`define TANH_LUT_2F38 16'h2F30
`define TANH_LUT_2F40 16'h2F38
`define TANH_LUT_2F48 16'h2F40
`define TANH_LUT_2F50 16'h2F48
`define TANH_LUT_2F58 16'h2F50
`define TANH_LUT_2F60 16'h2F58
`define TANH_LUT_2F68 16'h2F60
`define TANH_LUT_2F70 16'h2F67
`define TANH_LUT_2F78 16'h2F6F
`define TANH_LUT_2F80 16'h2F77
`define TANH_LUT_2F88 16'h2F7F
`define TANH_LUT_2F90 16'h2F87
`define TANH_LUT_2F98 16'h2F8F
`define TANH_LUT_2FA0 16'h2F97
`define TANH_LUT_2FA8 16'h2F9F
`define TANH_LUT_2FB0 16'h2FA7
`define TANH_LUT_2FB8 16'h2FAE
`define TANH_LUT_2FC0 16'h2FB6
`define TANH_LUT_2FC8 16'h2FBE
`define TANH_LUT_2FD0 16'h2FC6
`define TANH_LUT_2FD8 16'h2FCE
`define TANH_LUT_2FE0 16'h2FD6
`define TANH_LUT_2FE8 16'h2FDE
`define TANH_LUT_2FF0 16'h2FE6
`define TANH_LUT_2FF8 16'h2FEE
`define TANH_LUT_3000 16'h2FF5
`define TANH_LUT_3008 16'h3003
`define TANH_LUT_3010 16'h300A
`define TANH_LUT_3018 16'h3012
`define TANH_LUT_3020 16'h301A
`define TANH_LUT_3028 16'h3022
`define TANH_LUT_3030 16'h302A
`define TANH_LUT_3038 16'h3032
`define TANH_LUT_3040 16'h303A
`define TANH_LUT_3048 16'h3042
`define TANH_LUT_3050 16'h3049
`define TANH_LUT_3058 16'h3051
`define TANH_LUT_3060 16'h3059
`define TANH_LUT_3068 16'h3061
`define TANH_LUT_3070 16'h3069
`define TANH_LUT_3078 16'h3071
`define TANH_LUT_3080 16'h3078
`define TANH_LUT_3088 16'h3080
`define TANH_LUT_3090 16'h3088
`define TANH_LUT_3098 16'h3090
`define TANH_LUT_30A0 16'h3098
`define TANH_LUT_30A8 16'h30A0
`define TANH_LUT_30B0 16'h30A7
`define TANH_LUT_30B8 16'h30AF
`define TANH_LUT_30C0 16'h30B7
`define TANH_LUT_30C8 16'h30BF
`define TANH_LUT_30D0 16'h30C7
`define TANH_LUT_30D8 16'h30CF
`define TANH_LUT_30E0 16'h30D6
`define TANH_LUT_30E8 16'h30DE
`define TANH_LUT_30F0 16'h30E6
`define TANH_LUT_30F8 16'h30EE
`define TANH_LUT_3100 16'h30F6
`define TANH_LUT_3108 16'h30FD
`define TANH_LUT_3110 16'h3105
`define TANH_LUT_3118 16'h310D
`define TANH_LUT_3120 16'h3115
`define TANH_LUT_3128 16'h311D
`define TANH_LUT_3130 16'h3124
`define TANH_LUT_3138 16'h312C
`define TANH_LUT_3140 16'h3134
`define TANH_LUT_3148 16'h313C
`define TANH_LUT_3150 16'h3144
`define TANH_LUT_3158 16'h314B
`define TANH_LUT_3160 16'h3153
`define TANH_LUT_3168 16'h315B
`define TANH_LUT_3170 16'h3163
`define TANH_LUT_3178 16'h316B
`define TANH_LUT_3180 16'h3172
`define TANH_LUT_3188 16'h317A
`define TANH_LUT_3190 16'h3182
`define TANH_LUT_3198 16'h318A
`define TANH_LUT_31A0 16'h3191
`define TANH_LUT_31A8 16'h3199
`define TANH_LUT_31B0 16'h31A1
`define TANH_LUT_31B8 16'h31A9
`define TANH_LUT_31C0 16'h31B0
`define TANH_LUT_31C8 16'h31B8
`define TANH_LUT_31D0 16'h31C0
`define TANH_LUT_31D8 16'h31C8
`define TANH_LUT_31E0 16'h31CF
`define TANH_LUT_31E8 16'h31D7
`define TANH_LUT_31F0 16'h31DF
`define TANH_LUT_31F8 16'h31E7
`define TANH_LUT_3200 16'h31EE
`define TANH_LUT_3208 16'h31F6
`define TANH_LUT_3210 16'h31FE
`define TANH_LUT_3218 16'h3205
`define TANH_LUT_3220 16'h320D
`define TANH_LUT_3228 16'h3215
`define TANH_LUT_3230 16'h321D
`define TANH_LUT_3238 16'h3224
`define TANH_LUT_3240 16'h322C
`define TANH_LUT_3248 16'h3234
`define TANH_LUT_3250 16'h323B
`define TANH_LUT_3258 16'h3243
`define TANH_LUT_3260 16'h324B
`define TANH_LUT_3268 16'h3252
`define TANH_LUT_3270 16'h325A
`define TANH_LUT_3278 16'h3262
`define TANH_LUT_3280 16'h3269
`define TANH_LUT_3288 16'h3271
`define TANH_LUT_3290 16'h3279
`define TANH_LUT_3298 16'h3281
`define TANH_LUT_32A0 16'h3288
`define TANH_LUT_32A8 16'h3290
`define TANH_LUT_32B0 16'h3298
`define TANH_LUT_32B8 16'h329F
`define TANH_LUT_32C0 16'h32A7
`define TANH_LUT_32C8 16'h32AE
`define TANH_LUT_32D0 16'h32B6
`define TANH_LUT_32D8 16'h32BE
`define TANH_LUT_32E0 16'h32C5
`define TANH_LUT_32E8 16'h32CD
`define TANH_LUT_32F0 16'h32D5
`define TANH_LUT_32F8 16'h32DC
`define TANH_LUT_3300 16'h32E4
`define TANH_LUT_3308 16'h32EC
`define TANH_LUT_3310 16'h32F3
`define TANH_LUT_3318 16'h32FB
`define TANH_LUT_3320 16'h3302
`define TANH_LUT_3328 16'h330A
`define TANH_LUT_3330 16'h3312
`define TANH_LUT_3338 16'h3319
`define TANH_LUT_3340 16'h3321
`define TANH_LUT_3348 16'h3328
`define TANH_LUT_3350 16'h3330
`define TANH_LUT_3358 16'h3338
`define TANH_LUT_3360 16'h333F
`define TANH_LUT_3368 16'h3347
`define TANH_LUT_3370 16'h334E
`define TANH_LUT_3378 16'h3356
`define TANH_LUT_3380 16'h335E
`define TANH_LUT_3388 16'h3365
`define TANH_LUT_3390 16'h336D
`define TANH_LUT_3398 16'h3374
`define TANH_LUT_33A0 16'h337C
`define TANH_LUT_33A8 16'h3383
`define TANH_LUT_33B0 16'h338B
`define TANH_LUT_33B8 16'h3393
`define TANH_LUT_33C0 16'h339A
`define TANH_LUT_33C8 16'h33A2
`define TANH_LUT_33D0 16'h33A9
`define TANH_LUT_33D8 16'h33B1
`define TANH_LUT_33E0 16'h33B8
`define TANH_LUT_33E8 16'h33C0
`define TANH_LUT_33F0 16'h33C7
`define TANH_LUT_33F8 16'h33CF
`define TANH_LUT_3400 16'h33D6
`define TANH_LUT_3408 16'h33E5
`define TANH_LUT_3410 16'h33F4
`define TANH_LUT_3418 16'h3402
`define TANH_LUT_3420 16'h3409
`define TANH_LUT_3428 16'h3411
`define TANH_LUT_3430 16'h3418
`define TANH_LUT_3438 16'h3420
`define TANH_LUT_3440 16'h3427
`define TANH_LUT_3448 16'h342F
`define TANH_LUT_3450 16'h3436
`define TANH_LUT_3458 16'h343D
`define TANH_LUT_3460 16'h3445
`define TANH_LUT_3468 16'h344C
`define TANH_LUT_3470 16'h3454
`define TANH_LUT_3478 16'h345B
`define TANH_LUT_3480 16'h3463
`define TANH_LUT_3488 16'h346A
`define TANH_LUT_3490 16'h3471
`define TANH_LUT_3498 16'h3479
`define TANH_LUT_34A0 16'h3480
`define TANH_LUT_34A8 16'h3487
`define TANH_LUT_34B0 16'h348F
`define TANH_LUT_34B8 16'h3496
`define TANH_LUT_34C0 16'h349D
`define TANH_LUT_34C8 16'h34A5
`define TANH_LUT_34D0 16'h34AC
`define TANH_LUT_34D8 16'h34B3
`define TANH_LUT_34E0 16'h34BB
`define TANH_LUT_34E8 16'h34C2
`define TANH_LUT_34F0 16'h34C9
`define TANH_LUT_34F8 16'h34D1
`define TANH_LUT_3500 16'h34D8
`define TANH_LUT_3508 16'h34DF
`define TANH_LUT_3510 16'h34E6
`define TANH_LUT_3518 16'h34EE
`define TANH_LUT_3520 16'h34F5
`define TANH_LUT_3528 16'h34FC
`define TANH_LUT_3530 16'h3503
`define TANH_LUT_3538 16'h350B
`define TANH_LUT_3540 16'h3512
`define TANH_LUT_3548 16'h3519
`define TANH_LUT_3550 16'h3520
`define TANH_LUT_3558 16'h3527
`define TANH_LUT_3560 16'h352E
`define TANH_LUT_3568 16'h3536
`define TANH_LUT_3570 16'h353D
`define TANH_LUT_3578 16'h3544
`define TANH_LUT_3580 16'h354B
`define TANH_LUT_3588 16'h3552
`define TANH_LUT_3590 16'h3559
`define TANH_LUT_3598 16'h3560
`define TANH_LUT_35A0 16'h3567
`define TANH_LUT_35A8 16'h356F
`define TANH_LUT_35B0 16'h3576
`define TANH_LUT_35B8 16'h357D
`define TANH_LUT_35C0 16'h3584
`define TANH_LUT_35C8 16'h358B
`define TANH_LUT_35D0 16'h3592
`define TANH_LUT_35D8 16'h3599
`define TANH_LUT_35E0 16'h35A0
`define TANH_LUT_35E8 16'h35A7
`define TANH_LUT_35F0 16'h35AE
`define TANH_LUT_35F8 16'h35B5
`define TANH_LUT_3600 16'h35BC
`define TANH_LUT_3608 16'h35C3
`define TANH_LUT_3610 16'h35CA
`define TANH_LUT_3618 16'h35D1
`define TANH_LUT_3620 16'h35D8
`define TANH_LUT_3628 16'h35DF
`define TANH_LUT_3630 16'h35E5
`define TANH_LUT_3638 16'h35EC
`define TANH_LUT_3640 16'h35F3
`define TANH_LUT_3648 16'h35FA
`define TANH_LUT_3650 16'h3601
`define TANH_LUT_3658 16'h3608
`define TANH_LUT_3660 16'h360F
`define TANH_LUT_3668 16'h3616
`define TANH_LUT_3670 16'h361C
`define TANH_LUT_3678 16'h3623
`define TANH_LUT_3680 16'h362A
`define TANH_LUT_3688 16'h3631
`define TANH_LUT_3690 16'h3638
`define TANH_LUT_3698 16'h363F
`define TANH_LUT_36A0 16'h3645
`define TANH_LUT_36A8 16'h364C
`define TANH_LUT_36B0 16'h3653
`define TANH_LUT_36B8 16'h365A
`define TANH_LUT_36C0 16'h3660
`define TANH_LUT_36C8 16'h3667
`define TANH_LUT_36D0 16'h366E
`define TANH_LUT_36D8 16'h3674
`define TANH_LUT_36E0 16'h367B
`define TANH_LUT_36E8 16'h3682
`define TANH_LUT_36F0 16'h3688
`define TANH_LUT_36F8 16'h368F
`define TANH_LUT_3700 16'h3696
`define TANH_LUT_3708 16'h369C
`define TANH_LUT_3710 16'h36A3
`define TANH_LUT_3718 16'h36AA
`define TANH_LUT_3720 16'h36B0
`define TANH_LUT_3728 16'h36B7
`define TANH_LUT_3730 16'h36BD
`define TANH_LUT_3738 16'h36C4
`define TANH_LUT_3740 16'h36CB
`define TANH_LUT_3748 16'h36D1
`define TANH_LUT_3750 16'h36D8
`define TANH_LUT_3758 16'h36DE
`define TANH_LUT_3760 16'h36E5
`define TANH_LUT_3768 16'h36EB
`define TANH_LUT_3770 16'h36F2
`define TANH_LUT_3778 16'h36F8
`define TANH_LUT_3780 16'h36FF
`define TANH_LUT_3788 16'h3705
`define TANH_LUT_3790 16'h370C
`define TANH_LUT_3798 16'h3712
`define TANH_LUT_37A0 16'h3719
`define TANH_LUT_37A8 16'h371F
`define TANH_LUT_37B0 16'h3725
`define TANH_LUT_37B8 16'h372C
`define TANH_LUT_37C0 16'h3732
`define TANH_LUT_37C8 16'h3739
`define TANH_LUT_37D0 16'h373F
`define TANH_LUT_37D8 16'h3745
`define TANH_LUT_37E0 16'h374C
`define TANH_LUT_37E8 16'h3752
`define TANH_LUT_37F0 16'h3758
`define TANH_LUT_37F8 16'h375F
`define TANH_LUT_3800 16'h3765
`define TANH_LUT_3808 16'h3771
`define TANH_LUT_3810 16'h377E
`define TANH_LUT_3818 16'h378A
`define TANH_LUT_3820 16'h3797
`define TANH_LUT_3828 16'h37A3
`define TANH_LUT_3830 16'h37B0
`define TANH_LUT_3838 16'h37BC
`define TANH_LUT_3840 16'h37C8
`define TANH_LUT_3848 16'h37D4
`define TANH_LUT_3850 16'h37E0
`define TANH_LUT_3858 16'h37EC
`define TANH_LUT_3860 16'h37F9
`define TANH_LUT_3868 16'h3802
`define TANH_LUT_3870 16'h3808
`define TANH_LUT_3878 16'h380E
`define TANH_LUT_3880 16'h3814
`define TANH_LUT_3888 16'h381A
`define TANH_LUT_3890 16'h3820
`define TANH_LUT_3898 16'h3826
`define TANH_LUT_38A0 16'h382C
`define TANH_LUT_38A8 16'h3831
`define TANH_LUT_38B0 16'h3837
`define TANH_LUT_38B8 16'h383D
`define TANH_LUT_38C0 16'h3843
`define TANH_LUT_38C8 16'h3848
`define TANH_LUT_38D0 16'h384E
`define TANH_LUT_38D8 16'h3854
`define TANH_LUT_38E0 16'h3859
`define TANH_LUT_38E8 16'h385F
`define TANH_LUT_38F0 16'h3865
`define TANH_LUT_38F8 16'h386A
`define TANH_LUT_3900 16'h3870
`define TANH_LUT_3908 16'h3875
`define TANH_LUT_3910 16'h387B
`define TANH_LUT_3918 16'h3880
`define TANH_LUT_3920 16'h3886
`define TANH_LUT_3928 16'h388B
`define TANH_LUT_3930 16'h3891
`define TANH_LUT_3938 16'h3896
`define TANH_LUT_3940 16'h389B
`define TANH_LUT_3948 16'h38A1
`define TANH_LUT_3950 16'h38A6
`define TANH_LUT_3958 16'h38AB
`define TANH_LUT_3960 16'h38B1
`define TANH_LUT_3968 16'h38B6
`define TANH_LUT_3970 16'h38BB
`define TANH_LUT_3978 16'h38C0
`define TANH_LUT_3980 16'h38C5
`define TANH_LUT_3988 16'h38CB
`define TANH_LUT_3990 16'h38D0
`define TANH_LUT_3998 16'h38D5
`define TANH_LUT_39A0 16'h38DA
`define TANH_LUT_39A8 16'h38DF
`define TANH_LUT_39B0 16'h38E4
`define TANH_LUT_39B8 16'h38E9
`define TANH_LUT_39C0 16'h38EE
`define TANH_LUT_39C8 16'h38F3
`define TANH_LUT_39D0 16'h38F8
`define TANH_LUT_39D8 16'h38FD
`define TANH_LUT_39E0 16'h3902
`define TANH_LUT_39E8 16'h3906
`define TANH_LUT_39F0 16'h390B
`define TANH_LUT_39F8 16'h3910
`define TANH_LUT_3A00 16'h3915
`define TANH_LUT_3A08 16'h391A
`define TANH_LUT_3A10 16'h391E
`define TANH_LUT_3A18 16'h3923
`define TANH_LUT_3A20 16'h3928
`define TANH_LUT_3A28 16'h392C
`define TANH_LUT_3A30 16'h3931
`define TANH_LUT_3A38 16'h3936
`define TANH_LUT_3A40 16'h393A
`define TANH_LUT_3A48 16'h393F
`define TANH_LUT_3A50 16'h3943
`define TANH_LUT_3A58 16'h3948
`define TANH_LUT_3A60 16'h394C
`define TANH_LUT_3A68 16'h3951
`define TANH_LUT_3A70 16'h3955
`define TANH_LUT_3A78 16'h395A
`define TANH_LUT_3A80 16'h395E
`define TANH_LUT_3A88 16'h3963
`define TANH_LUT_3A90 16'h3967
`define TANH_LUT_3A98 16'h396B
`define TANH_LUT_3AA0 16'h3970
`define TANH_LUT_3AA8 16'h3974
`define TANH_LUT_3AB0 16'h3978
`define TANH_LUT_3AB8 16'h397C
`define TANH_LUT_3AC0 16'h3981
`define TANH_LUT_3AC8 16'h3985
`define TANH_LUT_3AD0 16'h3989
`define TANH_LUT_3AD8 16'h398D
`define TANH_LUT_3AE0 16'h3991
`define TANH_LUT_3AE8 16'h3995
`define TANH_LUT_3AF0 16'h3999
`define TANH_LUT_3AF8 16'h399E
`define TANH_LUT_3B00 16'h39A2
`define TANH_LUT_3B08 16'h39A6
`define TANH_LUT_3B10 16'h39AA
`define TANH_LUT_3B18 16'h39AE
`define TANH_LUT_3B20 16'h39B2
`define TANH_LUT_3B28 16'h39B6
`define TANH_LUT_3B30 16'h39B9
`define TANH_LUT_3B38 16'h39BD
`define TANH_LUT_3B40 16'h39C1
`define TANH_LUT_3B48 16'h39C5
`define TANH_LUT_3B50 16'h39C9
`define TANH_LUT_3B58 16'h39CD
`define TANH_LUT_3B60 16'h39D0
`define TANH_LUT_3B68 16'h39D4
`define TANH_LUT_3B70 16'h39D8
`define TANH_LUT_3B78 16'h39DC
`define TANH_LUT_3B80 16'h39DF
`define TANH_LUT_3B88 16'h39E3
`define TANH_LUT_3B90 16'h39E7
`define TANH_LUT_3B98 16'h39EA
`define TANH_LUT_3BA0 16'h39EE
`define TANH_LUT_3BA8 16'h39F2
`define TANH_LUT_3BB0 16'h39F5
`define TANH_LUT_3BB8 16'h39F9
`define TANH_LUT_3BC0 16'h39FC
`define TANH_LUT_3BC8 16'h3A00
`define TANH_LUT_3BD0 16'h3A03
`define TANH_LUT_3BD8 16'h3A07
`define TANH_LUT_3BE0 16'h3A0A
`define TANH_LUT_3BE8 16'h3A0E
`define TANH_LUT_3BF0 16'h3A11
`define TANH_LUT_3BF8 16'h3A14
`define TANH_LUT_3C00 16'h3A18
`define TANH_LUT_3C08 16'h3A1E
`define TANH_LUT_3C10 16'h3A25
`define TANH_LUT_3C18 16'h3A2C
`define TANH_LUT_3C20 16'h3A32
`define TANH_LUT_3C28 16'h3A38
`define TANH_LUT_3C30 16'h3A3F
`define TANH_LUT_3C38 16'h3A45
`define TANH_LUT_3C40 16'h3A4B
`define TANH_LUT_3C48 16'h3A51
`define TANH_LUT_3C50 16'h3A57
`define TANH_LUT_3C58 16'h3A5D
`define TANH_LUT_3C60 16'h3A63
`define TANH_LUT_3C68 16'h3A69
`define TANH_LUT_3C70 16'h3A6E
`define TANH_LUT_3C78 16'h3A74
`define TANH_LUT_3C80 16'h3A79
`define TANH_LUT_3C88 16'h3A7F
`define TANH_LUT_3C90 16'h3A84
`define TANH_LUT_3C98 16'h3A8A
`define TANH_LUT_3CA0 16'h3A8F
`define TANH_LUT_3CA8 16'h3A94
`define TANH_LUT_3CB0 16'h3A99
`define TANH_LUT_3CB8 16'h3A9E
`define TANH_LUT_3CC0 16'h3AA3
`define TANH_LUT_3CC8 16'h3AA8
`define TANH_LUT_3CD0 16'h3AAD
`define TANH_LUT_3CD8 16'h3AB2
`define TANH_LUT_3CE0 16'h3AB7
`define TANH_LUT_3CE8 16'h3ABC
`define TANH_LUT_3CF0 16'h3AC0
`define TANH_LUT_3CF8 16'h3AC5
`define TANH_LUT_3D00 16'h3AC9
`define TANH_LUT_3D08 16'h3ACE
`define TANH_LUT_3D10 16'h3AD2
`define TANH_LUT_3D18 16'h3AD6
`define TANH_LUT_3D20 16'h3ADB
`define TANH_LUT_3D28 16'h3ADF
`define TANH_LUT_3D30 16'h3AE3
`define TANH_LUT_3D38 16'h3AE7
`define TANH_LUT_3D40 16'h3AEB
`define TANH_LUT_3D48 16'h3AEF
`define TANH_LUT_3D50 16'h3AF3
`define TANH_LUT_3D58 16'h3AF7
`define TANH_LUT_3D60 16'h3AFB
`define TANH_LUT_3D68 16'h3AFF
`define TANH_LUT_3D70 16'h3B03
`define TANH_LUT_3D78 16'h3B06
`define TANH_LUT_3D80 16'h3B0A
`define TANH_LUT_3D88 16'h3B0D
`define TANH_LUT_3D90 16'h3B11
`define TANH_LUT_3D98 16'h3B15
`define TANH_LUT_3DA0 16'h3B18
`define TANH_LUT_3DA8 16'h3B1B
`define TANH_LUT_3DB0 16'h3B1F
`define TANH_LUT_3DB8 16'h3B22
`define TANH_LUT_3DC0 16'h3B25
`define TANH_LUT_3DC8 16'h3B28
`define TANH_LUT_3DD0 16'h3B2C
`define TANH_LUT_3DD8 16'h3B2F
`define TANH_LUT_3DE0 16'h3B32
`define TANH_LUT_3DE8 16'h3B35
`define TANH_LUT_3DF0 16'h3B38
`define TANH_LUT_3DF8 16'h3B3B
`define TANH_LUT_3E00 16'h3B3E
`define TANH_LUT_3E08 16'h3B41
`define TANH_LUT_3E10 16'h3B43
`define TANH_LUT_3E18 16'h3B46
`define TANH_LUT_3E20 16'h3B49
`define TANH_LUT_3E28 16'h3B4C
`define TANH_LUT_3E30 16'h3B4E
`define TANH_LUT_3E38 16'h3B51
`define TANH_LUT_3E40 16'h3B54
`define TANH_LUT_3E48 16'h3B56
`define TANH_LUT_3E50 16'h3B59
`define TANH_LUT_3E58 16'h3B5B
`define TANH_LUT_3E60 16'h3B5E
`define TANH_LUT_3E68 16'h3B60
`define TANH_LUT_3E70 16'h3B62
`define TANH_LUT_3E78 16'h3B65
`define TANH_LUT_3E80 16'h3B67
`define TANH_LUT_3E88 16'h3B69
`define TANH_LUT_3E90 16'h3B6C
`define TANH_LUT_3E98 16'h3B6E
`define TANH_LUT_3EA0 16'h3B70
`define TANH_LUT_3EA8 16'h3B72
`define TANH_LUT_3EB0 16'h3B74
`define TANH_LUT_3EB8 16'h3B76
`define TANH_LUT_3EC0 16'h3B78
`define TANH_LUT_3EC8 16'h3B7B
`define TANH_LUT_3ED0 16'h3B7D
`define TANH_LUT_3ED8 16'h3B7E
`define TANH_LUT_3EE0 16'h3B80
`define TANH_LUT_3EE8 16'h3B82
`define TANH_LUT_3EF0 16'h3B84
`define TANH_LUT_3EF8 16'h3B86
`define TANH_LUT_3F00 16'h3B88
`define TANH_LUT_3F08 16'h3B8A
`define TANH_LUT_3F10 16'h3B8C
`define TANH_LUT_3F18 16'h3B8D
`define TANH_LUT_3F20 16'h3B8F
`define TANH_LUT_3F28 16'h3B91
`define TANH_LUT_3F30 16'h3B92
`define TANH_LUT_3F38 16'h3B94
`define TANH_LUT_3F40 16'h3B96
`define TANH_LUT_3F48 16'h3B97
`define TANH_LUT_3F50 16'h3B99
`define TANH_LUT_3F58 16'h3B9A
`define TANH_LUT_3F60 16'h3B9C
`define TANH_LUT_3F68 16'h3B9D
`define TANH_LUT_3F70 16'h3B9F
`define TANH_LUT_3F78 16'h3BA0
`define TANH_LUT_3F80 16'h3BA2
`define TANH_LUT_3F88 16'h3BA3
`define TANH_LUT_3F90 16'h3BA5
`define TANH_LUT_3F98 16'h3BA6
`define TANH_LUT_3FA0 16'h3BA7
`define TANH_LUT_3FA8 16'h3BA9
`define TANH_LUT_3FB0 16'h3BAA
`define TANH_LUT_3FB8 16'h3BAB
`define TANH_LUT_3FC0 16'h3BAD
`define TANH_LUT_3FC8 16'h3BAE
`define TANH_LUT_3FD0 16'h3BAF
`define TANH_LUT_3FD8 16'h3BB0
`define TANH_LUT_3FE0 16'h3BB2
`define TANH_LUT_3FE8 16'h3BB3
`define TANH_LUT_3FF0 16'h3BB4
`define TANH_LUT_3FF8 16'h3BB5
`define TANH_LUT_4000 16'h3BB6
`define TANH_LUT_4008 16'h3BB9
`define TANH_LUT_4010 16'h3BBB
`define TANH_LUT_4018 16'h3BBD
`define TANH_LUT_4020 16'h3BBF
`define TANH_LUT_4028 16'h3BC1
`define TANH_LUT_4030 16'h3BC3
`define TANH_LUT_4038 16'h3BC5
`define TANH_LUT_4040 16'h3BC6
`define TANH_LUT_4048 16'h3BC8
`define TANH_LUT_4050 16'h3BCA
`define TANH_LUT_4058 16'h3BCB
`define TANH_LUT_4060 16'h3BCD
`define TANH_LUT_4068 16'h3BCF
`define TANH_LUT_4070 16'h3BD0
`define TANH_LUT_4078 16'h3BD2
`define TANH_LUT_4080 16'h3BD3
`define TANH_LUT_4088 16'h3BD4
`define TANH_LUT_4090 16'h3BD6
`define TANH_LUT_4098 16'h3BD7
`define TANH_LUT_40A0 16'h3BD8
`define TANH_LUT_40A8 16'h3BD9
`define TANH_LUT_40B0 16'h3BDB
`define TANH_LUT_40B8 16'h3BDC
`define TANH_LUT_40C0 16'h3BDD
`define TANH_LUT_40C8 16'h3BDE
`define TANH_LUT_40D0 16'h3BDF
`define TANH_LUT_40D8 16'h3BE0
`define TANH_LUT_40E0 16'h3BE1
`define TANH_LUT_40E8 16'h3BE2
`define TANH_LUT_40F0 16'h3BE3
`define TANH_LUT_40F8 16'h3BE4
`define TANH_LUT_4100 16'h3BE5
`define TANH_LUT_4108 16'h3BE5
`define TANH_LUT_4110 16'h3BE6
`define TANH_LUT_4118 16'h3BE7
`define TANH_LUT_4120 16'h3BE8
`define TANH_LUT_4128 16'h3BE9
`define TANH_LUT_4130 16'h3BE9
`define TANH_LUT_4138 16'h3BEA
`define TANH_LUT_4140 16'h3BEB
`define TANH_LUT_4148 16'h3BEB
`define TANH_LUT_4150 16'h3BEC
`define TANH_LUT_4158 16'h3BED
`define TANH_LUT_4160 16'h3BED
`define TANH_LUT_4168 16'h3BEE
`define TANH_LUT_4170 16'h3BEE
`define TANH_LUT_4178 16'h3BEF
`define TANH_LUT_4180 16'h3BEF
`define TANH_LUT_4188 16'h3BF0
`define TANH_LUT_4190 16'h3BF0
`define TANH_LUT_4198 16'h3BF1
`define TANH_LUT_41A0 16'h3BF1
`define TANH_LUT_41A8 16'h3BF2
`define TANH_LUT_41B0 16'h3BF2
`define TANH_LUT_41B8 16'h3BF3
`define TANH_LUT_41C0 16'h3BF3
`define TANH_LUT_41C8 16'h3BF3
`define TANH_LUT_41D0 16'h3BF4
`define TANH_LUT_41D8 16'h3BF4
`define TANH_LUT_41E0 16'h3BF5
`define TANH_LUT_41E8 16'h3BF5
`define TANH_LUT_41F0 16'h3BF5
`define TANH_LUT_41F8 16'h3BF6
`define TANH_LUT_4200 16'h3BF6
`define TANH_LUT_4208 16'h3BF6
`define TANH_LUT_4210 16'h3BF6
`define TANH_LUT_4218 16'h3BF7
`define TANH_LUT_4220 16'h3BF7
`define TANH_LUT_4228 16'h3BF7
`define TANH_LUT_4230 16'h3BF8
`define TANH_LUT_4238 16'h3BF8
`define TANH_LUT_4240 16'h3BF8
`define TANH_LUT_4248 16'h3BF8
`define TANH_LUT_4250 16'h3BF9
`define TANH_LUT_4258 16'h3BF9
`define TANH_LUT_4260 16'h3BF9
`define TANH_LUT_4268 16'h3BF9
`define TANH_LUT_4270 16'h3BF9
`define TANH_LUT_4278 16'h3BFA
`define TANH_LUT_4280 16'h3BFA
`define TANH_LUT_4288 16'h3BFA
`define TANH_LUT_4290 16'h3BFA
`define TANH_LUT_4298 16'h3BFA
`define TANH_LUT_42A0 16'h3BFB
`define TANH_LUT_42A8 16'h3BFB
`define TANH_LUT_42B0 16'h3BFB
`define TANH_LUT_42B8 16'h3BFB
`define TANH_LUT_42C0 16'h3BFB
`define TANH_LUT_42C8 16'h3BFB
`define TANH_LUT_42D0 16'h3BFB
`define TANH_LUT_42D8 16'h3BFC
`define TANH_LUT_8000 16'h8000
`define TANH_LUT_8008 16'h8008
`define TANH_LUT_8010 16'h8010
`define TANH_LUT_8018 16'h8018
`define TANH_LUT_8020 16'h8020
`define TANH_LUT_8028 16'h8028
`define TANH_LUT_8030 16'h8030
`define TANH_LUT_8038 16'h8038
`define TANH_LUT_8040 16'h8040
`define TANH_LUT_8048 16'h8048
`define TANH_LUT_8050 16'h8050
`define TANH_LUT_8058 16'h8058
`define TANH_LUT_8060 16'h8060
`define TANH_LUT_8068 16'h8068
`define TANH_LUT_8070 16'h8070
`define TANH_LUT_8078 16'h8078
`define TANH_LUT_8080 16'h8080
`define TANH_LUT_8088 16'h8088
`define TANH_LUT_8090 16'h8090
`define TANH_LUT_8098 16'h8098
`define TANH_LUT_80A0 16'h80A0
`define TANH_LUT_80A8 16'h80A8
`define TANH_LUT_80B0 16'h80B0
`define TANH_LUT_80B8 16'h80B8
`define TANH_LUT_80C0 16'h80C0
`define TANH_LUT_80C8 16'h80C8
`define TANH_LUT_80D0 16'h80D0
`define TANH_LUT_80D8 16'h80D8
`define TANH_LUT_80E0 16'h80E0
`define TANH_LUT_80E8 16'h80E8
`define TANH_LUT_80F0 16'h80F0
`define TANH_LUT_80F8 16'h80F8
`define TANH_LUT_8100 16'h8100
`define TANH_LUT_8108 16'h8108
`define TANH_LUT_8110 16'h8110
`define TANH_LUT_8118 16'h8118
`define TANH_LUT_8120 16'h8120
`define TANH_LUT_8128 16'h8128
`define TANH_LUT_8130 16'h8130
`define TANH_LUT_8138 16'h8138
`define TANH_LUT_8140 16'h8140
`define TANH_LUT_8148 16'h8148
`define TANH_LUT_8150 16'h8150
`define TANH_LUT_8158 16'h8158
`define TANH_LUT_8160 16'h8160
`define TANH_LUT_8168 16'h8168
`define TANH_LUT_8170 16'h8170
`define TANH_LUT_8178 16'h8178
`define TANH_LUT_8180 16'h8180
`define TANH_LUT_8188 16'h8188
`define TANH_LUT_8190 16'h8190
`define TANH_LUT_8198 16'h8198
`define TANH_LUT_81A0 16'h81A0
`define TANH_LUT_81A8 16'h81A8
`define TANH_LUT_81B0 16'h81B0
`define TANH_LUT_81B8 16'h81B8
`define TANH_LUT_81C0 16'h81C0
`define TANH_LUT_81C8 16'h81C8
`define TANH_LUT_81D0 16'h81D0
`define TANH_LUT_81D8 16'h81D8
`define TANH_LUT_81E0 16'h81E0
`define TANH_LUT_81E8 16'h81E8
`define TANH_LUT_81F0 16'h81F0
`define TANH_LUT_81F8 16'h81F8
`define TANH_LUT_8200 16'h8200
`define TANH_LUT_8208 16'h8208
`define TANH_LUT_8210 16'h8210
`define TANH_LUT_8218 16'h8218
`define TANH_LUT_8220 16'h8220
`define TANH_LUT_8228 16'h8228
`define TANH_LUT_8230 16'h8230
`define TANH_LUT_8238 16'h8238
`define TANH_LUT_8240 16'h8240
`define TANH_LUT_8248 16'h8248
`define TANH_LUT_8250 16'h8250
`define TANH_LUT_8258 16'h8258
`define TANH_LUT_8260 16'h8260
`define TANH_LUT_8268 16'h8268
`define TANH_LUT_8270 16'h8270
`define TANH_LUT_8278 16'h8278
`define TANH_LUT_8280 16'h8280
`define TANH_LUT_8288 16'h8288
`define TANH_LUT_8290 16'h8290
`define TANH_LUT_8298 16'h8298
`define TANH_LUT_82A0 16'h82A0
`define TANH_LUT_82A8 16'h82A8
`define TANH_LUT_82B0 16'h82B0
`define TANH_LUT_82B8 16'h82B8
`define TANH_LUT_82C0 16'h82C0
`define TANH_LUT_82C8 16'h82C8
`define TANH_LUT_82D0 16'h82D0
`define TANH_LUT_82D8 16'h82D8
`define TANH_LUT_82E0 16'h82E0
`define TANH_LUT_82E8 16'h82E8
`define TANH_LUT_82F0 16'h82F0
`define TANH_LUT_82F8 16'h82F8
`define TANH_LUT_8300 16'h8300
`define TANH_LUT_8308 16'h8308
`define TANH_LUT_8310 16'h8310
`define TANH_LUT_8318 16'h8318
`define TANH_LUT_8320 16'h8320
`define TANH_LUT_8328 16'h8328
`define TANH_LUT_8330 16'h8330
`define TANH_LUT_8338 16'h8338
`define TANH_LUT_8340 16'h8340
`define TANH_LUT_8348 16'h8348
`define TANH_LUT_8350 16'h8350
`define TANH_LUT_8358 16'h8358
`define TANH_LUT_8360 16'h8360
`define TANH_LUT_8368 16'h8368
`define TANH_LUT_8370 16'h8370
`define TANH_LUT_8378 16'h8378
`define TANH_LUT_8380 16'h8380
`define TANH_LUT_8388 16'h8388
`define TANH_LUT_8390 16'h8390
`define TANH_LUT_8398 16'h8398
`define TANH_LUT_83A0 16'h83A0
`define TANH_LUT_83A8 16'h83A8
`define TANH_LUT_83B0 16'h83B0
`define TANH_LUT_83B8 16'h83B8
`define TANH_LUT_83C0 16'h83C0
`define TANH_LUT_83C8 16'h83C8
`define TANH_LUT_83D0 16'h83D0
`define TANH_LUT_83D8 16'h83D8
`define TANH_LUT_83E0 16'h83E0
`define TANH_LUT_83E8 16'h83E8
`define TANH_LUT_83F0 16'h83F0
`define TANH_LUT_83F8 16'h83F8
`define TANH_LUT_8400 16'h8400
`define TANH_LUT_8408 16'h8408
`define TANH_LUT_8410 16'h8410
`define TANH_LUT_8418 16'h8418
`define TANH_LUT_8420 16'h8420
`define TANH_LUT_8428 16'h8428
`define TANH_LUT_8430 16'h8430
`define TANH_LUT_8438 16'h8438
`define TANH_LUT_8440 16'h8440
`define TANH_LUT_8448 16'h8448
`define TANH_LUT_8450 16'h8450
`define TANH_LUT_8458 16'h8458
`define TANH_LUT_8460 16'h8460
`define TANH_LUT_8468 16'h8468
`define TANH_LUT_8470 16'h8470
`define TANH_LUT_8478 16'h8478
`define TANH_LUT_8480 16'h8480
`define TANH_LUT_8488 16'h8488
`define TANH_LUT_8490 16'h8490
`define TANH_LUT_8498 16'h8498
`define TANH_LUT_84A0 16'h84A0
`define TANH_LUT_84A8 16'h84A8
`define TANH_LUT_84B0 16'h84B0
`define TANH_LUT_84B8 16'h84B8
`define TANH_LUT_84C0 16'h84C0
`define TANH_LUT_84C8 16'h84C8
`define TANH_LUT_84D0 16'h84D0
`define TANH_LUT_84D8 16'h84D8
`define TANH_LUT_84E0 16'h84E0
`define TANH_LUT_84E8 16'h84E8
`define TANH_LUT_84F0 16'h84F0
`define TANH_LUT_84F8 16'h84F8
`define TANH_LUT_8500 16'h8500
`define TANH_LUT_8508 16'h8508
`define TANH_LUT_8510 16'h8510
`define TANH_LUT_8518 16'h8518
`define TANH_LUT_8520 16'h8520
`define TANH_LUT_8528 16'h8528
`define TANH_LUT_8530 16'h8530
`define TANH_LUT_8538 16'h8538
`define TANH_LUT_8540 16'h8540
`define TANH_LUT_8548 16'h8548
`define TANH_LUT_8550 16'h8550
`define TANH_LUT_8558 16'h8558
`define TANH_LUT_8560 16'h8560
`define TANH_LUT_8568 16'h8568
`define TANH_LUT_8570 16'h8570
`define TANH_LUT_8578 16'h8578
`define TANH_LUT_8580 16'h8580
`define TANH_LUT_8588 16'h8588
`define TANH_LUT_8590 16'h8590
`define TANH_LUT_8598 16'h8598
`define TANH_LUT_85A0 16'h85A0
`define TANH_LUT_85A8 16'h85A8
`define TANH_LUT_85B0 16'h85B0
`define TANH_LUT_85B8 16'h85B8
`define TANH_LUT_85C0 16'h85C0
`define TANH_LUT_85C8 16'h85C8
`define TANH_LUT_85D0 16'h85D0
`define TANH_LUT_85D8 16'h85D8
`define TANH_LUT_85E0 16'h85E0
`define TANH_LUT_85E8 16'h85E8
`define TANH_LUT_85F0 16'h85F0
`define TANH_LUT_85F8 16'h85F8
`define TANH_LUT_8600 16'h8600
`define TANH_LUT_8608 16'h8608
`define TANH_LUT_8610 16'h8610
`define TANH_LUT_8618 16'h8618
`define TANH_LUT_8620 16'h8620
`define TANH_LUT_8628 16'h8628
`define TANH_LUT_8630 16'h8630
`define TANH_LUT_8638 16'h8638
`define TANH_LUT_8640 16'h8640
`define TANH_LUT_8648 16'h8648
`define TANH_LUT_8650 16'h8650
`define TANH_LUT_8658 16'h8658
`define TANH_LUT_8660 16'h8660
`define TANH_LUT_8668 16'h8668
`define TANH_LUT_8670 16'h8670
`define TANH_LUT_8678 16'h8678
`define TANH_LUT_8680 16'h8680
`define TANH_LUT_8688 16'h8688
`define TANH_LUT_8690 16'h8690
`define TANH_LUT_8698 16'h8698
`define TANH_LUT_86A0 16'h86A0
`define TANH_LUT_86A8 16'h86A8
`define TANH_LUT_86B0 16'h86B0
`define TANH_LUT_86B8 16'h86B8
`define TANH_LUT_86C0 16'h86C0
`define TANH_LUT_86C8 16'h86C8
`define TANH_LUT_86D0 16'h86D0
`define TANH_LUT_86D8 16'h86D8
`define TANH_LUT_86E0 16'h86E0
`define TANH_LUT_86E8 16'h86E8
`define TANH_LUT_86F0 16'h86F0
`define TANH_LUT_86F8 16'h86F8
`define TANH_LUT_8700 16'h8700
`define TANH_LUT_8708 16'h8708
`define TANH_LUT_8710 16'h8710
`define TANH_LUT_8718 16'h8718
`define TANH_LUT_8720 16'h8720
`define TANH_LUT_8728 16'h8728
`define TANH_LUT_8730 16'h8730
`define TANH_LUT_8738 16'h8738
`define TANH_LUT_8740 16'h8740
`define TANH_LUT_8748 16'h8748
`define TANH_LUT_8750 16'h8750
`define TANH_LUT_8758 16'h8758
`define TANH_LUT_8760 16'h8760
`define TANH_LUT_8768 16'h8768
`define TANH_LUT_8770 16'h8770
`define TANH_LUT_8778 16'h8778
`define TANH_LUT_8780 16'h8780
`define TANH_LUT_8788 16'h8788
`define TANH_LUT_8790 16'h8790
`define TANH_LUT_8798 16'h8798
`define TANH_LUT_87A0 16'h87A0
`define TANH_LUT_87A8 16'h87A8
`define TANH_LUT_87B0 16'h87B0
`define TANH_LUT_87B8 16'h87B8
`define TANH_LUT_87C0 16'h87C0
`define TANH_LUT_87C8 16'h87C8
`define TANH_LUT_87D0 16'h87D0
`define TANH_LUT_87D8 16'h87D8
`define TANH_LUT_87E0 16'h87E0
`define TANH_LUT_87E8 16'h87E8
`define TANH_LUT_87F0 16'h87F0
`define TANH_LUT_87F8 16'h87F8
`define TANH_LUT_8800 16'h8800
`define TANH_LUT_8808 16'h8808
`define TANH_LUT_8810 16'h8810
`define TANH_LUT_8818 16'h8818
`define TANH_LUT_8820 16'h8820
`define TANH_LUT_8828 16'h8828
`define TANH_LUT_8830 16'h8830
`define TANH_LUT_8838 16'h8838
`define TANH_LUT_8840 16'h8840
`define TANH_LUT_8848 16'h8848
`define TANH_LUT_8850 16'h8850
`define TANH_LUT_8858 16'h8858
`define TANH_LUT_8860 16'h8860
`define TANH_LUT_8868 16'h8868
`define TANH_LUT_8870 16'h8870
`define TANH_LUT_8878 16'h8878
`define TANH_LUT_8880 16'h8880
`define TANH_LUT_8888 16'h8888
`define TANH_LUT_8890 16'h8890
`define TANH_LUT_8898 16'h8898
`define TANH_LUT_88A0 16'h88A0
`define TANH_LUT_88A8 16'h88A8
`define TANH_LUT_88B0 16'h88B0
`define TANH_LUT_88B8 16'h88B8
`define TANH_LUT_88C0 16'h88C0
`define TANH_LUT_88C8 16'h88C8
`define TANH_LUT_88D0 16'h88D0
`define TANH_LUT_88D8 16'h88D8
`define TANH_LUT_88E0 16'h88E0
`define TANH_LUT_88E8 16'h88E8
`define TANH_LUT_88F0 16'h88F0
`define TANH_LUT_88F8 16'h88F8
`define TANH_LUT_8900 16'h8900
`define TANH_LUT_8908 16'h8908
`define TANH_LUT_8910 16'h8910
`define TANH_LUT_8918 16'h8918
`define TANH_LUT_8920 16'h8920
`define TANH_LUT_8928 16'h8928
`define TANH_LUT_8930 16'h8930
`define TANH_LUT_8938 16'h8938
`define TANH_LUT_8940 16'h8940
`define TANH_LUT_8948 16'h8948
`define TANH_LUT_8950 16'h8950
`define TANH_LUT_8958 16'h8958
`define TANH_LUT_8960 16'h8960
`define TANH_LUT_8968 16'h8968
`define TANH_LUT_8970 16'h8970
`define TANH_LUT_8978 16'h8978
`define TANH_LUT_8980 16'h8980
`define TANH_LUT_8988 16'h8988
`define TANH_LUT_8990 16'h8990
`define TANH_LUT_8998 16'h8998
`define TANH_LUT_89A0 16'h89A0
`define TANH_LUT_89A8 16'h89A8
`define TANH_LUT_89B0 16'h89B0
`define TANH_LUT_89B8 16'h89B8
`define TANH_LUT_89C0 16'h89C0
`define TANH_LUT_89C8 16'h89C8
`define TANH_LUT_89D0 16'h89D0
`define TANH_LUT_89D8 16'h89D8
`define TANH_LUT_89E0 16'h89E0
`define TANH_LUT_89E8 16'h89E8
`define TANH_LUT_89F0 16'h89F0
`define TANH_LUT_89F8 16'h89F8
`define TANH_LUT_8A00 16'h8A00
`define TANH_LUT_8A08 16'h8A08
`define TANH_LUT_8A10 16'h8A10
`define TANH_LUT_8A18 16'h8A18
`define TANH_LUT_8A20 16'h8A20
`define TANH_LUT_8A28 16'h8A28
`define TANH_LUT_8A30 16'h8A30
`define TANH_LUT_8A38 16'h8A38
`define TANH_LUT_8A40 16'h8A40
`define TANH_LUT_8A48 16'h8A48
`define TANH_LUT_8A50 16'h8A50
`define TANH_LUT_8A58 16'h8A58
`define TANH_LUT_8A60 16'h8A60
`define TANH_LUT_8A68 16'h8A68
`define TANH_LUT_8A70 16'h8A70
`define TANH_LUT_8A78 16'h8A78
`define TANH_LUT_8A80 16'h8A80
`define TANH_LUT_8A88 16'h8A88
`define TANH_LUT_8A90 16'h8A90
`define TANH_LUT_8A98 16'h8A98
`define TANH_LUT_8AA0 16'h8AA0
`define TANH_LUT_8AA8 16'h8AA8
`define TANH_LUT_8AB0 16'h8AB0
`define TANH_LUT_8AB8 16'h8AB8
`define TANH_LUT_8AC0 16'h8AC0
`define TANH_LUT_8AC8 16'h8AC8
`define TANH_LUT_8AD0 16'h8AD0
`define TANH_LUT_8AD8 16'h8AD8
`define TANH_LUT_8AE0 16'h8AE0
`define TANH_LUT_8AE8 16'h8AE8
`define TANH_LUT_8AF0 16'h8AF0
`define TANH_LUT_8AF8 16'h8AF8
`define TANH_LUT_8B00 16'h8B00
`define TANH_LUT_8B08 16'h8B08
`define TANH_LUT_8B10 16'h8B10
`define TANH_LUT_8B18 16'h8B18
`define TANH_LUT_8B20 16'h8B20
`define TANH_LUT_8B28 16'h8B28
`define TANH_LUT_8B30 16'h8B30
`define TANH_LUT_8B38 16'h8B38
`define TANH_LUT_8B40 16'h8B40
`define TANH_LUT_8B48 16'h8B48
`define TANH_LUT_8B50 16'h8B50
`define TANH_LUT_8B58 16'h8B58
`define TANH_LUT_8B60 16'h8B60
`define TANH_LUT_8B68 16'h8B68
`define TANH_LUT_8B70 16'h8B70
`define TANH_LUT_8B78 16'h8B78
`define TANH_LUT_8B80 16'h8B80
`define TANH_LUT_8B88 16'h8B88
`define TANH_LUT_8B90 16'h8B90
`define TANH_LUT_8B98 16'h8B98
`define TANH_LUT_8BA0 16'h8BA0
`define TANH_LUT_8BA8 16'h8BA8
`define TANH_LUT_8BB0 16'h8BB0
`define TANH_LUT_8BB8 16'h8BB8
`define TANH_LUT_8BC0 16'h8BC0
`define TANH_LUT_8BC8 16'h8BC8
`define TANH_LUT_8BD0 16'h8BD0
`define TANH_LUT_8BD8 16'h8BD8
`define TANH_LUT_8BE0 16'h8BE0
`define TANH_LUT_8BE8 16'h8BE8
`define TANH_LUT_8BF0 16'h8BF0
`define TANH_LUT_8BF8 16'h8BF8
`define TANH_LUT_8C00 16'h8C00
`define TANH_LUT_8C08 16'h8C08
`define TANH_LUT_8C10 16'h8C10
`define TANH_LUT_8C18 16'h8C18
`define TANH_LUT_8C20 16'h8C20
`define TANH_LUT_8C28 16'h8C28
`define TANH_LUT_8C30 16'h8C30
`define TANH_LUT_8C38 16'h8C38
`define TANH_LUT_8C40 16'h8C40
`define TANH_LUT_8C48 16'h8C48
`define TANH_LUT_8C50 16'h8C50
`define TANH_LUT_8C58 16'h8C58
`define TANH_LUT_8C60 16'h8C60
`define TANH_LUT_8C68 16'h8C68
`define TANH_LUT_8C70 16'h8C70
`define TANH_LUT_8C78 16'h8C78
`define TANH_LUT_8C80 16'h8C80
`define TANH_LUT_8C88 16'h8C88
`define TANH_LUT_8C90 16'h8C90
`define TANH_LUT_8C98 16'h8C98
`define TANH_LUT_8CA0 16'h8CA0
`define TANH_LUT_8CA8 16'h8CA8
`define TANH_LUT_8CB0 16'h8CB0
`define TANH_LUT_8CB8 16'h8CB8
`define TANH_LUT_8CC0 16'h8CC0
`define TANH_LUT_8CC8 16'h8CC8
`define TANH_LUT_8CD0 16'h8CD0
`define TANH_LUT_8CD8 16'h8CD8
`define TANH_LUT_8CE0 16'h8CE0
`define TANH_LUT_8CE8 16'h8CE8
`define TANH_LUT_8CF0 16'h8CF0
`define TANH_LUT_8CF8 16'h8CF8
`define TANH_LUT_8D00 16'h8D00
`define TANH_LUT_8D08 16'h8D08
`define TANH_LUT_8D10 16'h8D10
`define TANH_LUT_8D18 16'h8D18
`define TANH_LUT_8D20 16'h8D20
`define TANH_LUT_8D28 16'h8D28
`define TANH_LUT_8D30 16'h8D30
`define TANH_LUT_8D38 16'h8D38
`define TANH_LUT_8D40 16'h8D40
`define TANH_LUT_8D48 16'h8D48
`define TANH_LUT_8D50 16'h8D50
`define TANH_LUT_8D58 16'h8D58
`define TANH_LUT_8D60 16'h8D60
`define TANH_LUT_8D68 16'h8D68
`define TANH_LUT_8D70 16'h8D70
`define TANH_LUT_8D78 16'h8D78
`define TANH_LUT_8D80 16'h8D80
`define TANH_LUT_8D88 16'h8D88
`define TANH_LUT_8D90 16'h8D90
`define TANH_LUT_8D98 16'h8D98
`define TANH_LUT_8DA0 16'h8DA0
`define TANH_LUT_8DA8 16'h8DA8
`define TANH_LUT_8DB0 16'h8DB0
`define TANH_LUT_8DB8 16'h8DB8
`define TANH_LUT_8DC0 16'h8DC0
`define TANH_LUT_8DC8 16'h8DC8
`define TANH_LUT_8DD0 16'h8DD0
`define TANH_LUT_8DD8 16'h8DD8
`define TANH_LUT_8DE0 16'h8DE0
`define TANH_LUT_8DE8 16'h8DE8
`define TANH_LUT_8DF0 16'h8DF0
`define TANH_LUT_8DF8 16'h8DF8
`define TANH_LUT_8E00 16'h8E00
`define TANH_LUT_8E08 16'h8E08
`define TANH_LUT_8E10 16'h8E10
`define TANH_LUT_8E18 16'h8E18
`define TANH_LUT_8E20 16'h8E20
`define TANH_LUT_8E28 16'h8E28
`define TANH_LUT_8E30 16'h8E30
`define TANH_LUT_8E38 16'h8E38
`define TANH_LUT_8E40 16'h8E40
`define TANH_LUT_8E48 16'h8E48
`define TANH_LUT_8E50 16'h8E50
`define TANH_LUT_8E58 16'h8E58
`define TANH_LUT_8E60 16'h8E60
`define TANH_LUT_8E68 16'h8E68
`define TANH_LUT_8E70 16'h8E70
`define TANH_LUT_8E78 16'h8E78
`define TANH_LUT_8E80 16'h8E80
`define TANH_LUT_8E88 16'h8E88
`define TANH_LUT_8E90 16'h8E90
`define TANH_LUT_8E98 16'h8E98
`define TANH_LUT_8EA0 16'h8EA0
`define TANH_LUT_8EA8 16'h8EA8
`define TANH_LUT_8EB0 16'h8EB0
`define TANH_LUT_8EB8 16'h8EB8
`define TANH_LUT_8EC0 16'h8EC0
`define TANH_LUT_8EC8 16'h8EC8
`define TANH_LUT_8ED0 16'h8ED0
`define TANH_LUT_8ED8 16'h8ED8
`define TANH_LUT_8EE0 16'h8EE0
`define TANH_LUT_8EE8 16'h8EE8
`define TANH_LUT_8EF0 16'h8EF0
`define TANH_LUT_8EF8 16'h8EF8
`define TANH_LUT_8F00 16'h8F00
`define TANH_LUT_8F08 16'h8F08
`define TANH_LUT_8F10 16'h8F10
`define TANH_LUT_8F18 16'h8F18
`define TANH_LUT_8F20 16'h8F20
`define TANH_LUT_8F28 16'h8F28
`define TANH_LUT_8F30 16'h8F30
`define TANH_LUT_8F38 16'h8F38
`define TANH_LUT_8F40 16'h8F40
`define TANH_LUT_8F48 16'h8F48
`define TANH_LUT_8F50 16'h8F50
`define TANH_LUT_8F58 16'h8F58
`define TANH_LUT_8F60 16'h8F60
`define TANH_LUT_8F68 16'h8F68
`define TANH_LUT_8F70 16'h8F70
`define TANH_LUT_8F78 16'h8F78
`define TANH_LUT_8F80 16'h8F80
`define TANH_LUT_8F88 16'h8F88
`define TANH_LUT_8F90 16'h8F90
`define TANH_LUT_8F98 16'h8F98
`define TANH_LUT_8FA0 16'h8FA0
`define TANH_LUT_8FA8 16'h8FA8
`define TANH_LUT_8FB0 16'h8FB0
`define TANH_LUT_8FB8 16'h8FB8
`define TANH_LUT_8FC0 16'h8FC0
`define TANH_LUT_8FC8 16'h8FC8
`define TANH_LUT_8FD0 16'h8FD0
`define TANH_LUT_8FD8 16'h8FD8
`define TANH_LUT_8FE0 16'h8FE0
`define TANH_LUT_8FE8 16'h8FE8
`define TANH_LUT_8FF0 16'h8FF0
`define TANH_LUT_8FF8 16'h8FF8
`define TANH_LUT_9000 16'h9000
`define TANH_LUT_9008 16'h9008
`define TANH_LUT_9010 16'h9010
`define TANH_LUT_9018 16'h9018
`define TANH_LUT_9020 16'h9020
`define TANH_LUT_9028 16'h9028
`define TANH_LUT_9030 16'h9030
`define TANH_LUT_9038 16'h9038
`define TANH_LUT_9040 16'h9040
`define TANH_LUT_9048 16'h9048
`define TANH_LUT_9050 16'h9050
`define TANH_LUT_9058 16'h9058
`define TANH_LUT_9060 16'h9060
`define TANH_LUT_9068 16'h9068
`define TANH_LUT_9070 16'h9070
`define TANH_LUT_9078 16'h9078
`define TANH_LUT_9080 16'h9080
`define TANH_LUT_9088 16'h9088
`define TANH_LUT_9090 16'h9090
`define TANH_LUT_9098 16'h9098
`define TANH_LUT_90A0 16'h90A0
`define TANH_LUT_90A8 16'h90A8
`define TANH_LUT_90B0 16'h90B0
`define TANH_LUT_90B8 16'h90B8
`define TANH_LUT_90C0 16'h90C0
`define TANH_LUT_90C8 16'h90C8
`define TANH_LUT_90D0 16'h90D0
`define TANH_LUT_90D8 16'h90D8
`define TANH_LUT_90E0 16'h90E0
`define TANH_LUT_90E8 16'h90E8
`define TANH_LUT_90F0 16'h90F0
`define TANH_LUT_90F8 16'h90F8
`define TANH_LUT_9100 16'h9100
`define TANH_LUT_9108 16'h9108
`define TANH_LUT_9110 16'h9110
`define TANH_LUT_9118 16'h9118
`define TANH_LUT_9120 16'h9120
`define TANH_LUT_9128 16'h9128
`define TANH_LUT_9130 16'h9130
`define TANH_LUT_9138 16'h9138
`define TANH_LUT_9140 16'h9140
`define TANH_LUT_9148 16'h9148
`define TANH_LUT_9150 16'h9150
`define TANH_LUT_9158 16'h9158
`define TANH_LUT_9160 16'h9160
`define TANH_LUT_9168 16'h9168
`define TANH_LUT_9170 16'h9170
`define TANH_LUT_9178 16'h9178
`define TANH_LUT_9180 16'h9180
`define TANH_LUT_9188 16'h9188
`define TANH_LUT_9190 16'h9190
`define TANH_LUT_9198 16'h9198
`define TANH_LUT_91A0 16'h91A0
`define TANH_LUT_91A8 16'h91A8
`define TANH_LUT_91B0 16'h91B0
`define TANH_LUT_91B8 16'h91B8
`define TANH_LUT_91C0 16'h91C0
`define TANH_LUT_91C8 16'h91C8
`define TANH_LUT_91D0 16'h91D0
`define TANH_LUT_91D8 16'h91D8
`define TANH_LUT_91E0 16'h91E0
`define TANH_LUT_91E8 16'h91E8
`define TANH_LUT_91F0 16'h91F0
`define TANH_LUT_91F8 16'h91F8
`define TANH_LUT_9200 16'h9200
`define TANH_LUT_9208 16'h9208
`define TANH_LUT_9210 16'h9210
`define TANH_LUT_9218 16'h9218
`define TANH_LUT_9220 16'h9220
`define TANH_LUT_9228 16'h9228
`define TANH_LUT_9230 16'h9230
`define TANH_LUT_9238 16'h9238
`define TANH_LUT_9240 16'h9240
`define TANH_LUT_9248 16'h9248
`define TANH_LUT_9250 16'h9250
`define TANH_LUT_9258 16'h9258
`define TANH_LUT_9260 16'h9260
`define TANH_LUT_9268 16'h9268
`define TANH_LUT_9270 16'h9270
`define TANH_LUT_9278 16'h9278
`define TANH_LUT_9280 16'h9280
`define TANH_LUT_9288 16'h9288
`define TANH_LUT_9290 16'h9290
`define TANH_LUT_9298 16'h9298
`define TANH_LUT_92A0 16'h92A0
`define TANH_LUT_92A8 16'h92A8
`define TANH_LUT_92B0 16'h92B0
`define TANH_LUT_92B8 16'h92B8
`define TANH_LUT_92C0 16'h92C0
`define TANH_LUT_92C8 16'h92C8
`define TANH_LUT_92D0 16'h92D0
`define TANH_LUT_92D8 16'h92D8
`define TANH_LUT_92E0 16'h92E0
`define TANH_LUT_92E8 16'h92E8
`define TANH_LUT_92F0 16'h92F0
`define TANH_LUT_92F8 16'h92F8
`define TANH_LUT_9300 16'h9300
`define TANH_LUT_9308 16'h9308
`define TANH_LUT_9310 16'h9310
`define TANH_LUT_9318 16'h9318
`define TANH_LUT_9320 16'h9320
`define TANH_LUT_9328 16'h9328
`define TANH_LUT_9330 16'h9330
`define TANH_LUT_9338 16'h9338
`define TANH_LUT_9340 16'h9340
`define TANH_LUT_9348 16'h9348
`define TANH_LUT_9350 16'h9350
`define TANH_LUT_9358 16'h9358
`define TANH_LUT_9360 16'h9360
`define TANH_LUT_9368 16'h9368
`define TANH_LUT_9370 16'h9370
`define TANH_LUT_9378 16'h9378
`define TANH_LUT_9380 16'h9380
`define TANH_LUT_9388 16'h9388
`define TANH_LUT_9390 16'h9390
`define TANH_LUT_9398 16'h9398
`define TANH_LUT_93A0 16'h93A0
`define TANH_LUT_93A8 16'h93A8
`define TANH_LUT_93B0 16'h93B0
`define TANH_LUT_93B8 16'h93B8
`define TANH_LUT_93C0 16'h93C0
`define TANH_LUT_93C8 16'h93C8
`define TANH_LUT_93D0 16'h93D0
`define TANH_LUT_93D8 16'h93D8
`define TANH_LUT_93E0 16'h93E0
`define TANH_LUT_93E8 16'h93E8
`define TANH_LUT_93F0 16'h93F0
`define TANH_LUT_93F8 16'h93F8
`define TANH_LUT_9400 16'h9400
`define TANH_LUT_9408 16'h9408
`define TANH_LUT_9410 16'h9410
`define TANH_LUT_9418 16'h9418
`define TANH_LUT_9420 16'h9420
`define TANH_LUT_9428 16'h9428
`define TANH_LUT_9430 16'h9430
`define TANH_LUT_9438 16'h9438
`define TANH_LUT_9440 16'h9440
`define TANH_LUT_9448 16'h9448
`define TANH_LUT_9450 16'h9450
`define TANH_LUT_9458 16'h9458
`define TANH_LUT_9460 16'h9460
`define TANH_LUT_9468 16'h9468
`define TANH_LUT_9470 16'h9470
`define TANH_LUT_9478 16'h9478
`define TANH_LUT_9480 16'h9480
`define TANH_LUT_9488 16'h9488
`define TANH_LUT_9490 16'h9490
`define TANH_LUT_9498 16'h9498
`define TANH_LUT_94A0 16'h94A0
`define TANH_LUT_94A8 16'h94A8
`define TANH_LUT_94B0 16'h94B0
`define TANH_LUT_94B8 16'h94B8
`define TANH_LUT_94C0 16'h94C0
`define TANH_LUT_94C8 16'h94C8
`define TANH_LUT_94D0 16'h94D0
`define TANH_LUT_94D8 16'h94D8
`define TANH_LUT_94E0 16'h94E0
`define TANH_LUT_94E8 16'h94E8
`define TANH_LUT_94F0 16'h94F0
`define TANH_LUT_94F8 16'h94F8
`define TANH_LUT_9500 16'h9500
`define TANH_LUT_9508 16'h9508
`define TANH_LUT_9510 16'h9510
`define TANH_LUT_9518 16'h9518
`define TANH_LUT_9520 16'h9520
`define TANH_LUT_9528 16'h9528
`define TANH_LUT_9530 16'h9530
`define TANH_LUT_9538 16'h9538
`define TANH_LUT_9540 16'h9540
`define TANH_LUT_9548 16'h9548
`define TANH_LUT_9550 16'h9550
`define TANH_LUT_9558 16'h9558
`define TANH_LUT_9560 16'h9560
`define TANH_LUT_9568 16'h9568
`define TANH_LUT_9570 16'h9570
`define TANH_LUT_9578 16'h9578
`define TANH_LUT_9580 16'h9580
`define TANH_LUT_9588 16'h9588
`define TANH_LUT_9590 16'h9590
`define TANH_LUT_9598 16'h9598
`define TANH_LUT_95A0 16'h95A0
`define TANH_LUT_95A8 16'h95A8
`define TANH_LUT_95B0 16'h95B0
`define TANH_LUT_95B8 16'h95B8
`define TANH_LUT_95C0 16'h95C0
`define TANH_LUT_95C8 16'h95C8
`define TANH_LUT_95D0 16'h95D0
`define TANH_LUT_95D8 16'h95D8
`define TANH_LUT_95E0 16'h95E0
`define TANH_LUT_95E8 16'h95E8
`define TANH_LUT_95F0 16'h95F0
`define TANH_LUT_95F8 16'h95F8
`define TANH_LUT_9600 16'h9600
`define TANH_LUT_9608 16'h9608
`define TANH_LUT_9610 16'h9610
`define TANH_LUT_9618 16'h9618
`define TANH_LUT_9620 16'h9620
`define TANH_LUT_9628 16'h9628
`define TANH_LUT_9630 16'h9630
`define TANH_LUT_9638 16'h9638
`define TANH_LUT_9640 16'h9640
`define TANH_LUT_9648 16'h9648
`define TANH_LUT_9650 16'h9650
`define TANH_LUT_9658 16'h9658
`define TANH_LUT_9660 16'h9660
`define TANH_LUT_9668 16'h9668
`define TANH_LUT_9670 16'h9670
`define TANH_LUT_9678 16'h9678
`define TANH_LUT_9680 16'h9680
`define TANH_LUT_9688 16'h9688
`define TANH_LUT_9690 16'h9690
`define TANH_LUT_9698 16'h9698
`define TANH_LUT_96A0 16'h96A0
`define TANH_LUT_96A8 16'h96A8
`define TANH_LUT_96B0 16'h96B0
`define TANH_LUT_96B8 16'h96B8
`define TANH_LUT_96C0 16'h96C0
`define TANH_LUT_96C8 16'h96C8
`define TANH_LUT_96D0 16'h96D0
`define TANH_LUT_96D8 16'h96D8
`define TANH_LUT_96E0 16'h96E0
`define TANH_LUT_96E8 16'h96E8
`define TANH_LUT_96F0 16'h96F0
`define TANH_LUT_96F8 16'h96F8
`define TANH_LUT_9700 16'h9700
`define TANH_LUT_9708 16'h9708
`define TANH_LUT_9710 16'h9710
`define TANH_LUT_9718 16'h9718
`define TANH_LUT_9720 16'h9720
`define TANH_LUT_9728 16'h9728
`define TANH_LUT_9730 16'h9730
`define TANH_LUT_9738 16'h9738
`define TANH_LUT_9740 16'h9740
`define TANH_LUT_9748 16'h9748
`define TANH_LUT_9750 16'h9750
`define TANH_LUT_9758 16'h9758
`define TANH_LUT_9760 16'h9760
`define TANH_LUT_9768 16'h9768
`define TANH_LUT_9770 16'h9770
`define TANH_LUT_9778 16'h9778
`define TANH_LUT_9780 16'h9780
`define TANH_LUT_9788 16'h9788
`define TANH_LUT_9790 16'h9790
`define TANH_LUT_9798 16'h9798
`define TANH_LUT_97A0 16'h97A0
`define TANH_LUT_97A8 16'h97A8
`define TANH_LUT_97B0 16'h97B0
`define TANH_LUT_97B8 16'h97B8
`define TANH_LUT_97C0 16'h97C0
`define TANH_LUT_97C8 16'h97C8
`define TANH_LUT_97D0 16'h97D0
`define TANH_LUT_97D8 16'h97D8
`define TANH_LUT_97E0 16'h97E0
`define TANH_LUT_97E8 16'h97E8
`define TANH_LUT_97F0 16'h97F0
`define TANH_LUT_97F8 16'h97F8
`define TANH_LUT_9800 16'h9800
`define TANH_LUT_9808 16'h9808
`define TANH_LUT_9810 16'h9810
`define TANH_LUT_9818 16'h9818
`define TANH_LUT_9820 16'h9820
`define TANH_LUT_9828 16'h9828
`define TANH_LUT_9830 16'h9830
`define TANH_LUT_9838 16'h9838
`define TANH_LUT_9840 16'h9840
`define TANH_LUT_9848 16'h9848
`define TANH_LUT_9850 16'h9850
`define TANH_LUT_9858 16'h9858
`define TANH_LUT_9860 16'h9860
`define TANH_LUT_9868 16'h9868
`define TANH_LUT_9870 16'h9870
`define TANH_LUT_9878 16'h9878
`define TANH_LUT_9880 16'h9880
`define TANH_LUT_9888 16'h9888
`define TANH_LUT_9890 16'h9890
`define TANH_LUT_9898 16'h9898
`define TANH_LUT_98A0 16'h98A0
`define TANH_LUT_98A8 16'h98A8
`define TANH_LUT_98B0 16'h98B0
`define TANH_LUT_98B8 16'h98B8
`define TANH_LUT_98C0 16'h98C0
`define TANH_LUT_98C8 16'h98C8
`define TANH_LUT_98D0 16'h98D0
`define TANH_LUT_98D8 16'h98D8
`define TANH_LUT_98E0 16'h98E0
`define TANH_LUT_98E8 16'h98E8
`define TANH_LUT_98F0 16'h98F0
`define TANH_LUT_98F8 16'h98F8
`define TANH_LUT_9900 16'h9900
`define TANH_LUT_9908 16'h9908
`define TANH_LUT_9910 16'h9910
`define TANH_LUT_9918 16'h9918
`define TANH_LUT_9920 16'h9920
`define TANH_LUT_9928 16'h9928
`define TANH_LUT_9930 16'h9930
`define TANH_LUT_9938 16'h9938
`define TANH_LUT_9940 16'h9940
`define TANH_LUT_9948 16'h9948
`define TANH_LUT_9950 16'h9950
`define TANH_LUT_9958 16'h9958
`define TANH_LUT_9960 16'h9960
`define TANH_LUT_9968 16'h9968
`define TANH_LUT_9970 16'h9970
`define TANH_LUT_9978 16'h9978
`define TANH_LUT_9980 16'h9980
`define TANH_LUT_9988 16'h9988
`define TANH_LUT_9990 16'h9990
`define TANH_LUT_9998 16'h9998
`define TANH_LUT_99A0 16'h99A0
`define TANH_LUT_99A8 16'h99A8
`define TANH_LUT_99B0 16'h99B0
`define TANH_LUT_99B8 16'h99B8
`define TANH_LUT_99C0 16'h99C0
`define TANH_LUT_99C8 16'h99C8
`define TANH_LUT_99D0 16'h99D0
`define TANH_LUT_99D8 16'h99D8
`define TANH_LUT_99E0 16'h99E0
`define TANH_LUT_99E8 16'h99E8
`define TANH_LUT_99F0 16'h99F0
`define TANH_LUT_99F8 16'h99F8
`define TANH_LUT_9A00 16'h9A00
`define TANH_LUT_9A08 16'h9A08
`define TANH_LUT_9A10 16'h9A10
`define TANH_LUT_9A18 16'h9A18
`define TANH_LUT_9A20 16'h9A20
`define TANH_LUT_9A28 16'h9A28
`define TANH_LUT_9A30 16'h9A30
`define TANH_LUT_9A38 16'h9A38
`define TANH_LUT_9A40 16'h9A40
`define TANH_LUT_9A48 16'h9A48
`define TANH_LUT_9A50 16'h9A50
`define TANH_LUT_9A58 16'h9A58
`define TANH_LUT_9A60 16'h9A60
`define TANH_LUT_9A68 16'h9A68
`define TANH_LUT_9A70 16'h9A70
`define TANH_LUT_9A78 16'h9A78
`define TANH_LUT_9A80 16'h9A80
`define TANH_LUT_9A88 16'h9A88
`define TANH_LUT_9A90 16'h9A90
`define TANH_LUT_9A98 16'h9A98
`define TANH_LUT_9AA0 16'h9AA0
`define TANH_LUT_9AA8 16'h9AA8
`define TANH_LUT_9AB0 16'h9AB0
`define TANH_LUT_9AB8 16'h9AB8
`define TANH_LUT_9AC0 16'h9AC0
`define TANH_LUT_9AC8 16'h9AC8
`define TANH_LUT_9AD0 16'h9AD0
`define TANH_LUT_9AD8 16'h9AD8
`define TANH_LUT_9AE0 16'h9AE0
`define TANH_LUT_9AE8 16'h9AE8
`define TANH_LUT_9AF0 16'h9AF0
`define TANH_LUT_9AF8 16'h9AF8
`define TANH_LUT_9B00 16'h9B00
`define TANH_LUT_9B08 16'h9B08
`define TANH_LUT_9B10 16'h9B10
`define TANH_LUT_9B18 16'h9B18
`define TANH_LUT_9B20 16'h9B20
`define TANH_LUT_9B28 16'h9B28
`define TANH_LUT_9B30 16'h9B30
`define TANH_LUT_9B38 16'h9B38
`define TANH_LUT_9B40 16'h9B40
`define TANH_LUT_9B48 16'h9B48
`define TANH_LUT_9B50 16'h9B50
`define TANH_LUT_9B58 16'h9B58
`define TANH_LUT_9B60 16'h9B60
`define TANH_LUT_9B68 16'h9B68
`define TANH_LUT_9B70 16'h9B70
`define TANH_LUT_9B78 16'h9B78
`define TANH_LUT_9B80 16'h9B80
`define TANH_LUT_9B88 16'h9B88
`define TANH_LUT_9B90 16'h9B90
`define TANH_LUT_9B98 16'h9B98
`define TANH_LUT_9BA0 16'h9BA0
`define TANH_LUT_9BA8 16'h9BA8
`define TANH_LUT_9BB0 16'h9BB0
`define TANH_LUT_9BB8 16'h9BB8
`define TANH_LUT_9BC0 16'h9BC0
`define TANH_LUT_9BC8 16'h9BC8
`define TANH_LUT_9BD0 16'h9BD0
`define TANH_LUT_9BD8 16'h9BD8
`define TANH_LUT_9BE0 16'h9BE0
`define TANH_LUT_9BE8 16'h9BE8
`define TANH_LUT_9BF0 16'h9BF0
`define TANH_LUT_9BF8 16'h9BF8
`define TANH_LUT_9C00 16'h9C00
`define TANH_LUT_9C08 16'h9C08
`define TANH_LUT_9C10 16'h9C10
`define TANH_LUT_9C18 16'h9C18
`define TANH_LUT_9C20 16'h9C20
`define TANH_LUT_9C28 16'h9C28
`define TANH_LUT_9C30 16'h9C30
`define TANH_LUT_9C38 16'h9C38
`define TANH_LUT_9C40 16'h9C40
`define TANH_LUT_9C48 16'h9C48
`define TANH_LUT_9C50 16'h9C50
`define TANH_LUT_9C58 16'h9C58
`define TANH_LUT_9C60 16'h9C60
`define TANH_LUT_9C68 16'h9C68
`define TANH_LUT_9C70 16'h9C70
`define TANH_LUT_9C78 16'h9C78
`define TANH_LUT_9C80 16'h9C80
`define TANH_LUT_9C88 16'h9C88
`define TANH_LUT_9C90 16'h9C90
`define TANH_LUT_9C98 16'h9C98
`define TANH_LUT_9CA0 16'h9CA0
`define TANH_LUT_9CA8 16'h9CA8
`define TANH_LUT_9CB0 16'h9CB0
`define TANH_LUT_9CB8 16'h9CB8
`define TANH_LUT_9CC0 16'h9CC0
`define TANH_LUT_9CC8 16'h9CC8
`define TANH_LUT_9CD0 16'h9CD0
`define TANH_LUT_9CD8 16'h9CD8
`define TANH_LUT_9CE0 16'h9CE0
`define TANH_LUT_9CE8 16'h9CE8
`define TANH_LUT_9CF0 16'h9CF0
`define TANH_LUT_9CF8 16'h9CF8
`define TANH_LUT_9D00 16'h9D00
`define TANH_LUT_9D08 16'h9D08
`define TANH_LUT_9D10 16'h9D10
`define TANH_LUT_9D18 16'h9D18
`define TANH_LUT_9D20 16'h9D20
`define TANH_LUT_9D28 16'h9D28
`define TANH_LUT_9D30 16'h9D30
`define TANH_LUT_9D38 16'h9D38
`define TANH_LUT_9D40 16'h9D40
`define TANH_LUT_9D48 16'h9D48
`define TANH_LUT_9D50 16'h9D50
`define TANH_LUT_9D58 16'h9D58
`define TANH_LUT_9D60 16'h9D60
`define TANH_LUT_9D68 16'h9D68
`define TANH_LUT_9D70 16'h9D70
`define TANH_LUT_9D78 16'h9D78
`define TANH_LUT_9D80 16'h9D80
`define TANH_LUT_9D88 16'h9D88
`define TANH_LUT_9D90 16'h9D90
`define TANH_LUT_9D98 16'h9D98
`define TANH_LUT_9DA0 16'h9DA0
`define TANH_LUT_9DA8 16'h9DA8
`define TANH_LUT_9DB0 16'h9DB0
`define TANH_LUT_9DB8 16'h9DB8
`define TANH_LUT_9DC0 16'h9DC0
`define TANH_LUT_9DC8 16'h9DC8
`define TANH_LUT_9DD0 16'h9DD0
`define TANH_LUT_9DD8 16'h9DD8
`define TANH_LUT_9DE0 16'h9DE0
`define TANH_LUT_9DE8 16'h9DE8
`define TANH_LUT_9DF0 16'h9DF0
`define TANH_LUT_9DF8 16'h9DF8
`define TANH_LUT_9E00 16'h9E00
`define TANH_LUT_9E08 16'h9E08
`define TANH_LUT_9E10 16'h9E10
`define TANH_LUT_9E18 16'h9E18
`define TANH_LUT_9E20 16'h9E20
`define TANH_LUT_9E28 16'h9E28
`define TANH_LUT_9E30 16'h9E30
`define TANH_LUT_9E38 16'h9E38
`define TANH_LUT_9E40 16'h9E40
`define TANH_LUT_9E48 16'h9E48
`define TANH_LUT_9E50 16'h9E50
`define TANH_LUT_9E58 16'h9E58
`define TANH_LUT_9E60 16'h9E60
`define TANH_LUT_9E68 16'h9E68
`define TANH_LUT_9E70 16'h9E70
`define TANH_LUT_9E78 16'h9E78
`define TANH_LUT_9E80 16'h9E80
`define TANH_LUT_9E88 16'h9E88
`define TANH_LUT_9E90 16'h9E90
`define TANH_LUT_9E98 16'h9E98
`define TANH_LUT_9EA0 16'h9EA0
`define TANH_LUT_9EA8 16'h9EA8
`define TANH_LUT_9EB0 16'h9EB0
`define TANH_LUT_9EB8 16'h9EB8
`define TANH_LUT_9EC0 16'h9EC0
`define TANH_LUT_9EC8 16'h9EC8
`define TANH_LUT_9ED0 16'h9ED0
`define TANH_LUT_9ED8 16'h9ED8
`define TANH_LUT_9EE0 16'h9EE0
`define TANH_LUT_9EE8 16'h9EE8
`define TANH_LUT_9EF0 16'h9EF0
`define TANH_LUT_9EF8 16'h9EF8
`define TANH_LUT_9F00 16'h9F00
`define TANH_LUT_9F08 16'h9F08
`define TANH_LUT_9F10 16'h9F10
`define TANH_LUT_9F18 16'h9F18
`define TANH_LUT_9F20 16'h9F20
`define TANH_LUT_9F28 16'h9F28
`define TANH_LUT_9F30 16'h9F30
`define TANH_LUT_9F38 16'h9F38
`define TANH_LUT_9F40 16'h9F40
`define TANH_LUT_9F48 16'h9F48
`define TANH_LUT_9F50 16'h9F50
`define TANH_LUT_9F58 16'h9F58
`define TANH_LUT_9F60 16'h9F60
`define TANH_LUT_9F68 16'h9F68
`define TANH_LUT_9F70 16'h9F70
`define TANH_LUT_9F78 16'h9F78
`define TANH_LUT_9F80 16'h9F80
`define TANH_LUT_9F88 16'h9F88
`define TANH_LUT_9F90 16'h9F90
`define TANH_LUT_9F98 16'h9F98
`define TANH_LUT_9FA0 16'h9FA0
`define TANH_LUT_9FA8 16'h9FA8
`define TANH_LUT_9FB0 16'h9FB0
`define TANH_LUT_9FB8 16'h9FB8
`define TANH_LUT_9FC0 16'h9FC0
`define TANH_LUT_9FC8 16'h9FC8
`define TANH_LUT_9FD0 16'h9FD0
`define TANH_LUT_9FD8 16'h9FD8
`define TANH_LUT_9FE0 16'h9FE0
`define TANH_LUT_9FE8 16'h9FE8
`define TANH_LUT_9FF0 16'h9FF0
`define TANH_LUT_9FF8 16'h9FF8
`define TANH_LUT_A000 16'hA000
`define TANH_LUT_A008 16'hA008
`define TANH_LUT_A010 16'hA010
`define TANH_LUT_A018 16'hA018
`define TANH_LUT_A020 16'hA020
`define TANH_LUT_A028 16'hA028
`define TANH_LUT_A030 16'hA030
`define TANH_LUT_A038 16'hA038
`define TANH_LUT_A040 16'hA040
`define TANH_LUT_A048 16'hA048
`define TANH_LUT_A050 16'hA050
`define TANH_LUT_A058 16'hA058
`define TANH_LUT_A060 16'hA060
`define TANH_LUT_A068 16'hA068
`define TANH_LUT_A070 16'hA070
`define TANH_LUT_A078 16'hA078
`define TANH_LUT_A080 16'hA080
`define TANH_LUT_A088 16'hA088
`define TANH_LUT_A090 16'hA090
`define TANH_LUT_A098 16'hA098
`define TANH_LUT_A0A0 16'hA0A0
`define TANH_LUT_A0A8 16'hA0A8
`define TANH_LUT_A0B0 16'hA0B0
`define TANH_LUT_A0B8 16'hA0B8
`define TANH_LUT_A0C0 16'hA0C0
`define TANH_LUT_A0C8 16'hA0C8
`define TANH_LUT_A0D0 16'hA0D0
`define TANH_LUT_A0D8 16'hA0D8
`define TANH_LUT_A0E0 16'hA0E0
`define TANH_LUT_A0E8 16'hA0E8
`define TANH_LUT_A0F0 16'hA0F0
`define TANH_LUT_A0F8 16'hA0F8
`define TANH_LUT_A100 16'hA100
`define TANH_LUT_A108 16'hA108
`define TANH_LUT_A110 16'hA110
`define TANH_LUT_A118 16'hA118
`define TANH_LUT_A120 16'hA120
`define TANH_LUT_A128 16'hA128
`define TANH_LUT_A130 16'hA130
`define TANH_LUT_A138 16'hA138
`define TANH_LUT_A140 16'hA140
`define TANH_LUT_A148 16'hA148
`define TANH_LUT_A150 16'hA150
`define TANH_LUT_A158 16'hA158
`define TANH_LUT_A160 16'hA160
`define TANH_LUT_A168 16'hA168
`define TANH_LUT_A170 16'hA170
`define TANH_LUT_A178 16'hA178
`define TANH_LUT_A180 16'hA180
`define TANH_LUT_A188 16'hA188
`define TANH_LUT_A190 16'hA190
`define TANH_LUT_A198 16'hA198
`define TANH_LUT_A1A0 16'hA1A0
`define TANH_LUT_A1A8 16'hA1A8
`define TANH_LUT_A1B0 16'hA1B0
`define TANH_LUT_A1B8 16'hA1B8
`define TANH_LUT_A1C0 16'hA1C0
`define TANH_LUT_A1C8 16'hA1C8
`define TANH_LUT_A1D0 16'hA1D0
`define TANH_LUT_A1D8 16'hA1D8
`define TANH_LUT_A1E0 16'hA1E0
`define TANH_LUT_A1E8 16'hA1E8
`define TANH_LUT_A1F0 16'hA1F0
`define TANH_LUT_A1F8 16'hA1F8
`define TANH_LUT_A200 16'hA200
`define TANH_LUT_A208 16'hA208
`define TANH_LUT_A210 16'hA210
`define TANH_LUT_A218 16'hA218
`define TANH_LUT_A220 16'hA220
`define TANH_LUT_A228 16'hA228
`define TANH_LUT_A230 16'hA230
`define TANH_LUT_A238 16'hA238
`define TANH_LUT_A240 16'hA240
`define TANH_LUT_A248 16'hA248
`define TANH_LUT_A250 16'hA250
`define TANH_LUT_A258 16'hA258
`define TANH_LUT_A260 16'hA260
`define TANH_LUT_A268 16'hA268
`define TANH_LUT_A270 16'hA270
`define TANH_LUT_A278 16'hA278
`define TANH_LUT_A280 16'hA280
`define TANH_LUT_A288 16'hA288
`define TANH_LUT_A290 16'hA290
`define TANH_LUT_A298 16'hA298
`define TANH_LUT_A2A0 16'hA2A0
`define TANH_LUT_A2A8 16'hA2A8
`define TANH_LUT_A2B0 16'hA2B0
`define TANH_LUT_A2B8 16'hA2B8
`define TANH_LUT_A2C0 16'hA2C0
`define TANH_LUT_A2C8 16'hA2C8
`define TANH_LUT_A2D0 16'hA2D0
`define TANH_LUT_A2D8 16'hA2D8
`define TANH_LUT_A2E0 16'hA2E0
`define TANH_LUT_A2E8 16'hA2E8
`define TANH_LUT_A2F0 16'hA2F0
`define TANH_LUT_A2F8 16'hA2F8
`define TANH_LUT_A300 16'hA300
`define TANH_LUT_A308 16'hA308
`define TANH_LUT_A310 16'hA310
`define TANH_LUT_A318 16'hA318
`define TANH_LUT_A320 16'hA320
`define TANH_LUT_A328 16'hA328
`define TANH_LUT_A330 16'hA330
`define TANH_LUT_A338 16'hA338
`define TANH_LUT_A340 16'hA340
`define TANH_LUT_A348 16'hA348
`define TANH_LUT_A350 16'hA350
`define TANH_LUT_A358 16'hA358
`define TANH_LUT_A360 16'hA360
`define TANH_LUT_A368 16'hA368
`define TANH_LUT_A370 16'hA370
`define TANH_LUT_A378 16'hA378
`define TANH_LUT_A380 16'hA380
`define TANH_LUT_A388 16'hA388
`define TANH_LUT_A390 16'hA390
`define TANH_LUT_A398 16'hA398
`define TANH_LUT_A3A0 16'hA3A0
`define TANH_LUT_A3A8 16'hA3A8
`define TANH_LUT_A3B0 16'hA3B0
`define TANH_LUT_A3B8 16'hA3B8
`define TANH_LUT_A3C0 16'hA3C0
`define TANH_LUT_A3C8 16'hA3C8
`define TANH_LUT_A3D0 16'hA3D0
`define TANH_LUT_A3D8 16'hA3D8
`define TANH_LUT_A3E0 16'hA3E0
`define TANH_LUT_A3E8 16'hA3E8
`define TANH_LUT_A3F0 16'hA3F0
`define TANH_LUT_A3F8 16'hA3F8
`define TANH_LUT_A400 16'hA400
`define TANH_LUT_A408 16'hA408
`define TANH_LUT_A410 16'hA410
`define TANH_LUT_A418 16'hA418
`define TANH_LUT_A420 16'hA420
`define TANH_LUT_A428 16'hA428
`define TANH_LUT_A430 16'hA430
`define TANH_LUT_A438 16'hA438
`define TANH_LUT_A440 16'hA440
`define TANH_LUT_A448 16'hA448
`define TANH_LUT_A450 16'hA450
`define TANH_LUT_A458 16'hA458
`define TANH_LUT_A460 16'hA460
`define TANH_LUT_A468 16'hA468
`define TANH_LUT_A470 16'hA470
`define TANH_LUT_A478 16'hA478
`define TANH_LUT_A480 16'hA480
`define TANH_LUT_A488 16'hA488
`define TANH_LUT_A490 16'hA490
`define TANH_LUT_A498 16'hA498
`define TANH_LUT_A4A0 16'hA4A0
`define TANH_LUT_A4A8 16'hA4A8
`define TANH_LUT_A4B0 16'hA4B0
`define TANH_LUT_A4B8 16'hA4B8
`define TANH_LUT_A4C0 16'hA4C0
`define TANH_LUT_A4C8 16'hA4C8
`define TANH_LUT_A4D0 16'hA4D0
`define TANH_LUT_A4D8 16'hA4D8
`define TANH_LUT_A4E0 16'hA4E0
`define TANH_LUT_A4E8 16'hA4E8
`define TANH_LUT_A4F0 16'hA4F0
`define TANH_LUT_A4F8 16'hA4F8
`define TANH_LUT_A500 16'hA500
`define TANH_LUT_A508 16'hA508
`define TANH_LUT_A510 16'hA510
`define TANH_LUT_A518 16'hA518
`define TANH_LUT_A520 16'hA520
`define TANH_LUT_A528 16'hA528
`define TANH_LUT_A530 16'hA530
`define TANH_LUT_A538 16'hA538
`define TANH_LUT_A540 16'hA540
`define TANH_LUT_A548 16'hA548
`define TANH_LUT_A550 16'hA550
`define TANH_LUT_A558 16'hA558
`define TANH_LUT_A560 16'hA560
`define TANH_LUT_A568 16'hA568
`define TANH_LUT_A570 16'hA570
`define TANH_LUT_A578 16'hA578
`define TANH_LUT_A580 16'hA580
`define TANH_LUT_A588 16'hA588
`define TANH_LUT_A590 16'hA590
`define TANH_LUT_A598 16'hA598
`define TANH_LUT_A5A0 16'hA5A0
`define TANH_LUT_A5A8 16'hA5A8
`define TANH_LUT_A5B0 16'hA5B0
`define TANH_LUT_A5B8 16'hA5B8
`define TANH_LUT_A5C0 16'hA5C0
`define TANH_LUT_A5C8 16'hA5C8
`define TANH_LUT_A5D0 16'hA5D0
`define TANH_LUT_A5D8 16'hA5D8
`define TANH_LUT_A5E0 16'hA5E0
`define TANH_LUT_A5E8 16'hA5E8
`define TANH_LUT_A5F0 16'hA5F0
`define TANH_LUT_A5F8 16'hA5F8
`define TANH_LUT_A600 16'hA600
`define TANH_LUT_A608 16'hA608
`define TANH_LUT_A610 16'hA610
`define TANH_LUT_A618 16'hA618
`define TANH_LUT_A620 16'hA620
`define TANH_LUT_A628 16'hA628
`define TANH_LUT_A630 16'hA630
`define TANH_LUT_A638 16'hA638
`define TANH_LUT_A640 16'hA640
`define TANH_LUT_A648 16'hA648
`define TANH_LUT_A650 16'hA650
`define TANH_LUT_A658 16'hA658
`define TANH_LUT_A660 16'hA660
`define TANH_LUT_A668 16'hA668
`define TANH_LUT_A670 16'hA670
`define TANH_LUT_A678 16'hA678
`define TANH_LUT_A680 16'hA680
`define TANH_LUT_A688 16'hA688
`define TANH_LUT_A690 16'hA690
`define TANH_LUT_A698 16'hA698
`define TANH_LUT_A6A0 16'hA6A0
`define TANH_LUT_A6A8 16'hA6A8
`define TANH_LUT_A6B0 16'hA6B0
`define TANH_LUT_A6B8 16'hA6B8
`define TANH_LUT_A6C0 16'hA6C0
`define TANH_LUT_A6C8 16'hA6C8
`define TANH_LUT_A6D0 16'hA6D0
`define TANH_LUT_A6D8 16'hA6D8
`define TANH_LUT_A6E0 16'hA6E0
`define TANH_LUT_A6E8 16'hA6E8
`define TANH_LUT_A6F0 16'hA6F0
`define TANH_LUT_A6F8 16'hA6F8
`define TANH_LUT_A700 16'hA700
`define TANH_LUT_A708 16'hA708
`define TANH_LUT_A710 16'hA710
`define TANH_LUT_A718 16'hA718
`define TANH_LUT_A720 16'hA720
`define TANH_LUT_A728 16'hA728
`define TANH_LUT_A730 16'hA730
`define TANH_LUT_A738 16'hA738
`define TANH_LUT_A740 16'hA740
`define TANH_LUT_A748 16'hA747
`define TANH_LUT_A750 16'hA74F
`define TANH_LUT_A758 16'hA757
`define TANH_LUT_A760 16'hA75F
`define TANH_LUT_A768 16'hA767
`define TANH_LUT_A770 16'hA76F
`define TANH_LUT_A778 16'hA777
`define TANH_LUT_A780 16'hA77F
`define TANH_LUT_A788 16'hA787
`define TANH_LUT_A790 16'hA78F
`define TANH_LUT_A798 16'hA797
`define TANH_LUT_A7A0 16'hA79F
`define TANH_LUT_A7A8 16'hA7A7
`define TANH_LUT_A7B0 16'hA7AF
`define TANH_LUT_A7B8 16'hA7B7
`define TANH_LUT_A7C0 16'hA7BF
`define TANH_LUT_A7C8 16'hA7C7
`define TANH_LUT_A7D0 16'hA7CF
`define TANH_LUT_A7D8 16'hA7D7
`define TANH_LUT_A7E0 16'hA7DF
`define TANH_LUT_A7E8 16'hA7E7
`define TANH_LUT_A7F0 16'hA7EF
`define TANH_LUT_A7F8 16'hA7F7
`define TANH_LUT_A800 16'hA7FF
`define TANH_LUT_A808 16'hA808
`define TANH_LUT_A810 16'hA810
`define TANH_LUT_A818 16'hA818
`define TANH_LUT_A820 16'hA820
`define TANH_LUT_A828 16'hA828
`define TANH_LUT_A830 16'hA830
`define TANH_LUT_A838 16'hA838
`define TANH_LUT_A840 16'hA840
`define TANH_LUT_A848 16'hA848
`define TANH_LUT_A850 16'hA850
`define TANH_LUT_A858 16'hA858
`define TANH_LUT_A860 16'hA860
`define TANH_LUT_A868 16'hA868
`define TANH_LUT_A870 16'hA870
`define TANH_LUT_A878 16'hA878
`define TANH_LUT_A880 16'hA880
`define TANH_LUT_A888 16'hA888
`define TANH_LUT_A890 16'hA890
`define TANH_LUT_A898 16'hA897
`define TANH_LUT_A8A0 16'hA89F
`define TANH_LUT_A8A8 16'hA8A7
`define TANH_LUT_A8B0 16'hA8AF
`define TANH_LUT_A8B8 16'hA8B7
`define TANH_LUT_A8C0 16'hA8BF
`define TANH_LUT_A8C8 16'hA8C7
`define TANH_LUT_A8D0 16'hA8CF
`define TANH_LUT_A8D8 16'hA8D7
`define TANH_LUT_A8E0 16'hA8DF
`define TANH_LUT_A8E8 16'hA8E7
`define TANH_LUT_A8F0 16'hA8EF
`define TANH_LUT_A8F8 16'hA8F7
`define TANH_LUT_A900 16'hA8FF
`define TANH_LUT_A908 16'hA907
`define TANH_LUT_A910 16'hA90F
`define TANH_LUT_A918 16'hA917
`define TANH_LUT_A920 16'hA91F
`define TANH_LUT_A928 16'hA927
`define TANH_LUT_A930 16'hA92F
`define TANH_LUT_A938 16'hA937
`define TANH_LUT_A940 16'hA93F
`define TANH_LUT_A948 16'hA947
`define TANH_LUT_A950 16'hA94F
`define TANH_LUT_A958 16'hA957
`define TANH_LUT_A960 16'hA95F
`define TANH_LUT_A968 16'hA967
`define TANH_LUT_A970 16'hA96F
`define TANH_LUT_A978 16'hA977
`define TANH_LUT_A980 16'hA97F
`define TANH_LUT_A988 16'hA987
`define TANH_LUT_A990 16'hA98F
`define TANH_LUT_A998 16'hA997
`define TANH_LUT_A9A0 16'hA99F
`define TANH_LUT_A9A8 16'hA9A7
`define TANH_LUT_A9B0 16'hA9AF
`define TANH_LUT_A9B8 16'hA9B7
`define TANH_LUT_A9C0 16'hA9BF
`define TANH_LUT_A9C8 16'hA9C7
`define TANH_LUT_A9D0 16'hA9CF
`define TANH_LUT_A9D8 16'hA9D7
`define TANH_LUT_A9E0 16'hA9DF
`define TANH_LUT_A9E8 16'hA9E7
`define TANH_LUT_A9F0 16'hA9EF
`define TANH_LUT_A9F8 16'hA9F7
`define TANH_LUT_AA00 16'hA9FF
`define TANH_LUT_AA08 16'hAA07
`define TANH_LUT_AA10 16'hAA0F
`define TANH_LUT_AA18 16'hAA17
`define TANH_LUT_AA20 16'hAA1F
`define TANH_LUT_AA28 16'hAA27
`define TANH_LUT_AA30 16'hAA2F
`define TANH_LUT_AA38 16'hAA37
`define TANH_LUT_AA40 16'hAA3F
`define TANH_LUT_AA48 16'hAA47
`define TANH_LUT_AA50 16'hAA4F
`define TANH_LUT_AA58 16'hAA57
`define TANH_LUT_AA60 16'hAA5F
`define TANH_LUT_AA68 16'hAA67
`define TANH_LUT_AA70 16'hAA6F
`define TANH_LUT_AA78 16'hAA77
`define TANH_LUT_AA80 16'hAA7F
`define TANH_LUT_AA88 16'hAA87
`define TANH_LUT_AA90 16'hAA8F
`define TANH_LUT_AA98 16'hAA97
`define TANH_LUT_AAA0 16'hAA9E
`define TANH_LUT_AAA8 16'hAAA6
`define TANH_LUT_AAB0 16'hAAAE
`define TANH_LUT_AAB8 16'hAAB6
`define TANH_LUT_AAC0 16'hAABE
`define TANH_LUT_AAC8 16'hAAC6
`define TANH_LUT_AAD0 16'hAACE
`define TANH_LUT_AAD8 16'hAAD6
`define TANH_LUT_AAE0 16'hAADE
`define TANH_LUT_AAE8 16'hAAE6
`define TANH_LUT_AAF0 16'hAAEE
`define TANH_LUT_AAF8 16'hAAF6
`define TANH_LUT_AB00 16'hAAFE
`define TANH_LUT_AB08 16'hAB06
`define TANH_LUT_AB10 16'hAB0E
`define TANH_LUT_AB18 16'hAB16
`define TANH_LUT_AB20 16'hAB1E
`define TANH_LUT_AB28 16'hAB26
`define TANH_LUT_AB30 16'hAB2E
`define TANH_LUT_AB38 16'hAB36
`define TANH_LUT_AB40 16'hAB3E
`define TANH_LUT_AB48 16'hAB46
`define TANH_LUT_AB50 16'hAB4E
`define TANH_LUT_AB58 16'hAB56
`define TANH_LUT_AB60 16'hAB5E
`define TANH_LUT_AB68 16'hAB66
`define TANH_LUT_AB70 16'hAB6E
`define TANH_LUT_AB78 16'hAB76
`define TANH_LUT_AB80 16'hAB7E
`define TANH_LUT_AB88 16'hAB86
`define TANH_LUT_AB90 16'hAB8E
`define TANH_LUT_AB98 16'hAB96
`define TANH_LUT_ABA0 16'hAB9E
`define TANH_LUT_ABA8 16'hABA6
`define TANH_LUT_ABB0 16'hABAE
`define TANH_LUT_ABB8 16'hABB6
`define TANH_LUT_ABC0 16'hABBE
`define TANH_LUT_ABC8 16'hABC6
`define TANH_LUT_ABD0 16'hABCE
`define TANH_LUT_ABD8 16'hABD5
`define TANH_LUT_ABE0 16'hABDD
`define TANH_LUT_ABE8 16'hABE5
`define TANH_LUT_ABF0 16'hABED
`define TANH_LUT_ABF8 16'hABF5
`define TANH_LUT_AC00 16'hABFD
`define TANH_LUT_AC08 16'hAC07
`define TANH_LUT_AC10 16'hAC0F
`define TANH_LUT_AC18 16'hAC17
`define TANH_LUT_AC20 16'hAC1F
`define TANH_LUT_AC28 16'hAC27
`define TANH_LUT_AC30 16'hAC2E
`define TANH_LUT_AC38 16'hAC36
`define TANH_LUT_AC40 16'hAC3E
`define TANH_LUT_AC48 16'hAC46
`define TANH_LUT_AC50 16'hAC4E
`define TANH_LUT_AC58 16'hAC56
`define TANH_LUT_AC60 16'hAC5E
`define TANH_LUT_AC68 16'hAC66
`define TANH_LUT_AC70 16'hAC6E
`define TANH_LUT_AC78 16'hAC76
`define TANH_LUT_AC80 16'hAC7E
`define TANH_LUT_AC88 16'hAC86
`define TANH_LUT_AC90 16'hAC8E
`define TANH_LUT_AC98 16'hAC96
`define TANH_LUT_ACA0 16'hAC9E
`define TANH_LUT_ACA8 16'hACA6
`define TANH_LUT_ACB0 16'hACAE
`define TANH_LUT_ACB8 16'hACB6
`define TANH_LUT_ACC0 16'hACBE
`define TANH_LUT_ACC8 16'hACC6
`define TANH_LUT_ACD0 16'hACCE
`define TANH_LUT_ACD8 16'hACD6
`define TANH_LUT_ACE0 16'hACDE
`define TANH_LUT_ACE8 16'hACE6
`define TANH_LUT_ACF0 16'hACED
`define TANH_LUT_ACF8 16'hACF5
`define TANH_LUT_AD00 16'hACFD
`define TANH_LUT_AD08 16'hAD05
`define TANH_LUT_AD10 16'hAD0D
`define TANH_LUT_AD18 16'hAD15
`define TANH_LUT_AD20 16'hAD1D
`define TANH_LUT_AD28 16'hAD25
`define TANH_LUT_AD30 16'hAD2D
`define TANH_LUT_AD38 16'hAD35
`define TANH_LUT_AD40 16'hAD3D
`define TANH_LUT_AD48 16'hAD45
`define TANH_LUT_AD50 16'hAD4D
`define TANH_LUT_AD58 16'hAD55
`define TANH_LUT_AD60 16'hAD5D
`define TANH_LUT_AD68 16'hAD65
`define TANH_LUT_AD70 16'hAD6D
`define TANH_LUT_AD78 16'hAD75
`define TANH_LUT_AD80 16'hAD7D
`define TANH_LUT_AD88 16'hAD84
`define TANH_LUT_AD90 16'hAD8C
`define TANH_LUT_AD98 16'hAD94
`define TANH_LUT_ADA0 16'hAD9C
`define TANH_LUT_ADA8 16'hADA4
`define TANH_LUT_ADB0 16'hADAC
`define TANH_LUT_ADB8 16'hADB4
`define TANH_LUT_ADC0 16'hADBC
`define TANH_LUT_ADC8 16'hADC4
`define TANH_LUT_ADD0 16'hADCC
`define TANH_LUT_ADD8 16'hADD4
`define TANH_LUT_ADE0 16'hADDC
`define TANH_LUT_ADE8 16'hADE4
`define TANH_LUT_ADF0 16'hADEC
`define TANH_LUT_ADF8 16'hADF4
`define TANH_LUT_AE00 16'hADFC
`define TANH_LUT_AE08 16'hAE03
`define TANH_LUT_AE10 16'hAE0B
`define TANH_LUT_AE18 16'hAE13
`define TANH_LUT_AE20 16'hAE1B
`define TANH_LUT_AE28 16'hAE23
`define TANH_LUT_AE30 16'hAE2B
`define TANH_LUT_AE38 16'hAE33
`define TANH_LUT_AE40 16'hAE3B
`define TANH_LUT_AE48 16'hAE43
`define TANH_LUT_AE50 16'hAE4B
`define TANH_LUT_AE58 16'hAE53
`define TANH_LUT_AE60 16'hAE5B
`define TANH_LUT_AE68 16'hAE63
`define TANH_LUT_AE70 16'hAE6A
`define TANH_LUT_AE78 16'hAE72
`define TANH_LUT_AE80 16'hAE7A
`define TANH_LUT_AE88 16'hAE82
`define TANH_LUT_AE90 16'hAE8A
`define TANH_LUT_AE98 16'hAE92
`define TANH_LUT_AEA0 16'hAE9A
`define TANH_LUT_AEA8 16'hAEA2
`define TANH_LUT_AEB0 16'hAEAA
`define TANH_LUT_AEB8 16'hAEB2
`define TANH_LUT_AEC0 16'hAEBA
`define TANH_LUT_AEC8 16'hAEC2
`define TANH_LUT_AED0 16'hAEC9
`define TANH_LUT_AED8 16'hAED1
`define TANH_LUT_AEE0 16'hAED9
`define TANH_LUT_AEE8 16'hAEE1
`define TANH_LUT_AEF0 16'hAEE9
`define TANH_LUT_AEF8 16'hAEF1
`define TANH_LUT_AF00 16'hAEF9
`define TANH_LUT_AF08 16'hAF01
`define TANH_LUT_AF10 16'hAF09
`define TANH_LUT_AF18 16'hAF11
`define TANH_LUT_AF20 16'hAF19
`define TANH_LUT_AF28 16'hAF20
`define TANH_LUT_AF30 16'hAF28
`define TANH_LUT_AF38 16'hAF30
`define TANH_LUT_AF40 16'hAF38
`define TANH_LUT_AF48 16'hAF40
`define TANH_LUT_AF50 16'hAF48
`define TANH_LUT_AF58 16'hAF50
`define TANH_LUT_AF60 16'hAF58
`define TANH_LUT_AF68 16'hAF60
`define TANH_LUT_AF70 16'hAF67
`define TANH_LUT_AF78 16'hAF6F
`define TANH_LUT_AF80 16'hAF77
`define TANH_LUT_AF88 16'hAF7F
`define TANH_LUT_AF90 16'hAF87
`define TANH_LUT_AF98 16'hAF8F
`define TANH_LUT_AFA0 16'hAF97
`define TANH_LUT_AFA8 16'hAF9F
`define TANH_LUT_AFB0 16'hAFA7
`define TANH_LUT_AFB8 16'hAFAE
`define TANH_LUT_AFC0 16'hAFB6
`define TANH_LUT_AFC8 16'hAFBE
`define TANH_LUT_AFD0 16'hAFC6
`define TANH_LUT_AFD8 16'hAFCE
`define TANH_LUT_AFE0 16'hAFD6
`define TANH_LUT_AFE8 16'hAFDE
`define TANH_LUT_AFF0 16'hAFE6
`define TANH_LUT_AFF8 16'hAFEE
`define TANH_LUT_B000 16'hAFF5
`define TANH_LUT_B008 16'hB003
`define TANH_LUT_B010 16'hB00A
`define TANH_LUT_B018 16'hB012
`define TANH_LUT_B020 16'hB01A
`define TANH_LUT_B028 16'hB022
`define TANH_LUT_B030 16'hB02A
`define TANH_LUT_B038 16'hB032
`define TANH_LUT_B040 16'hB03A
`define TANH_LUT_B048 16'hB042
`define TANH_LUT_B050 16'hB049
`define TANH_LUT_B058 16'hB051
`define TANH_LUT_B060 16'hB059
`define TANH_LUT_B068 16'hB061
`define TANH_LUT_B070 16'hB069
`define TANH_LUT_B078 16'hB071
`define TANH_LUT_B080 16'hB078
`define TANH_LUT_B088 16'hB080
`define TANH_LUT_B090 16'hB088
`define TANH_LUT_B098 16'hB090
`define TANH_LUT_B0A0 16'hB098
`define TANH_LUT_B0A8 16'hB0A0
`define TANH_LUT_B0B0 16'hB0A7
`define TANH_LUT_B0B8 16'hB0AF
`define TANH_LUT_B0C0 16'hB0B7
`define TANH_LUT_B0C8 16'hB0BF
`define TANH_LUT_B0D0 16'hB0C7
`define TANH_LUT_B0D8 16'hB0CF
`define TANH_LUT_B0E0 16'hB0D6
`define TANH_LUT_B0E8 16'hB0DE
`define TANH_LUT_B0F0 16'hB0E6
`define TANH_LUT_B0F8 16'hB0EE
`define TANH_LUT_B100 16'hB0F6
`define TANH_LUT_B108 16'hB0FD
`define TANH_LUT_B110 16'hB105
`define TANH_LUT_B118 16'hB10D
`define TANH_LUT_B120 16'hB115
`define TANH_LUT_B128 16'hB11D
`define TANH_LUT_B130 16'hB124
`define TANH_LUT_B138 16'hB12C
`define TANH_LUT_B140 16'hB134
`define TANH_LUT_B148 16'hB13C
`define TANH_LUT_B150 16'hB144
`define TANH_LUT_B158 16'hB14B
`define TANH_LUT_B160 16'hB153
`define TANH_LUT_B168 16'hB15B
`define TANH_LUT_B170 16'hB163
`define TANH_LUT_B178 16'hB16B
`define TANH_LUT_B180 16'hB172
`define TANH_LUT_B188 16'hB17A
`define TANH_LUT_B190 16'hB182
`define TANH_LUT_B198 16'hB18A
`define TANH_LUT_B1A0 16'hB191
`define TANH_LUT_B1A8 16'hB199
`define TANH_LUT_B1B0 16'hB1A1
`define TANH_LUT_B1B8 16'hB1A9
`define TANH_LUT_B1C0 16'hB1B0
`define TANH_LUT_B1C8 16'hB1B8
`define TANH_LUT_B1D0 16'hB1C0
`define TANH_LUT_B1D8 16'hB1C8
`define TANH_LUT_B1E0 16'hB1CF
`define TANH_LUT_B1E8 16'hB1D7
`define TANH_LUT_B1F0 16'hB1DF
`define TANH_LUT_B1F8 16'hB1E7
`define TANH_LUT_B200 16'hB1EE
`define TANH_LUT_B208 16'hB1F6
`define TANH_LUT_B210 16'hB1FE
`define TANH_LUT_B218 16'hB205
`define TANH_LUT_B220 16'hB20D
`define TANH_LUT_B228 16'hB215
`define TANH_LUT_B230 16'hB21D
`define TANH_LUT_B238 16'hB224
`define TANH_LUT_B240 16'hB22C
`define TANH_LUT_B248 16'hB234
`define TANH_LUT_B250 16'hB23B
`define TANH_LUT_B258 16'hB243
`define TANH_LUT_B260 16'hB24B
`define TANH_LUT_B268 16'hB252
`define TANH_LUT_B270 16'hB25A
`define TANH_LUT_B278 16'hB262
`define TANH_LUT_B280 16'hB269
`define TANH_LUT_B288 16'hB271
`define TANH_LUT_B290 16'hB279
`define TANH_LUT_B298 16'hB281
`define TANH_LUT_B2A0 16'hB288
`define TANH_LUT_B2A8 16'hB290
`define TANH_LUT_B2B0 16'hB298
`define TANH_LUT_B2B8 16'hB29F
`define TANH_LUT_B2C0 16'hB2A7
`define TANH_LUT_B2C8 16'hB2AE
`define TANH_LUT_B2D0 16'hB2B6
`define TANH_LUT_B2D8 16'hB2BE
`define TANH_LUT_B2E0 16'hB2C5
`define TANH_LUT_B2E8 16'hB2CD
`define TANH_LUT_B2F0 16'hB2D5
`define TANH_LUT_B2F8 16'hB2DC
`define TANH_LUT_B300 16'hB2E4
`define TANH_LUT_B308 16'hB2EC
`define TANH_LUT_B310 16'hB2F3
`define TANH_LUT_B318 16'hB2FB
`define TANH_LUT_B320 16'hB302
`define TANH_LUT_B328 16'hB30A
`define TANH_LUT_B330 16'hB312
`define TANH_LUT_B338 16'hB319
`define TANH_LUT_B340 16'hB321
`define TANH_LUT_B348 16'hB328
`define TANH_LUT_B350 16'hB330
`define TANH_LUT_B358 16'hB338
`define TANH_LUT_B360 16'hB33F
`define TANH_LUT_B368 16'hB347
`define TANH_LUT_B370 16'hB34E
`define TANH_LUT_B378 16'hB356
`define TANH_LUT_B380 16'hB35E
`define TANH_LUT_B388 16'hB365
`define TANH_LUT_B390 16'hB36D
`define TANH_LUT_B398 16'hB374
`define TANH_LUT_B3A0 16'hB37C
`define TANH_LUT_B3A8 16'hB383
`define TANH_LUT_B3B0 16'hB38B
`define TANH_LUT_B3B8 16'hB393
`define TANH_LUT_B3C0 16'hB39A
`define TANH_LUT_B3C8 16'hB3A2
`define TANH_LUT_B3D0 16'hB3A9
`define TANH_LUT_B3D8 16'hB3B1
`define TANH_LUT_B3E0 16'hB3B8
`define TANH_LUT_B3E8 16'hB3C0
`define TANH_LUT_B3F0 16'hB3C7
`define TANH_LUT_B3F8 16'hB3CF
`define TANH_LUT_B400 16'hB3D6
`define TANH_LUT_B408 16'hB3E5
`define TANH_LUT_B410 16'hB3F4
`define TANH_LUT_B418 16'hB402
`define TANH_LUT_B420 16'hB409
`define TANH_LUT_B428 16'hB411
`define TANH_LUT_B430 16'hB418
`define TANH_LUT_B438 16'hB420
`define TANH_LUT_B440 16'hB427
`define TANH_LUT_B448 16'hB42F
`define TANH_LUT_B450 16'hB436
`define TANH_LUT_B458 16'hB43D
`define TANH_LUT_B460 16'hB445
`define TANH_LUT_B468 16'hB44C
`define TANH_LUT_B470 16'hB454
`define TANH_LUT_B478 16'hB45B
`define TANH_LUT_B480 16'hB463
`define TANH_LUT_B488 16'hB46A
`define TANH_LUT_B490 16'hB471
`define TANH_LUT_B498 16'hB479
`define TANH_LUT_B4A0 16'hB480
`define TANH_LUT_B4A8 16'hB487
`define TANH_LUT_B4B0 16'hB48F
`define TANH_LUT_B4B8 16'hB496
`define TANH_LUT_B4C0 16'hB49D
`define TANH_LUT_B4C8 16'hB4A5
`define TANH_LUT_B4D0 16'hB4AC
`define TANH_LUT_B4D8 16'hB4B3
`define TANH_LUT_B4E0 16'hB4BB
`define TANH_LUT_B4E8 16'hB4C2
`define TANH_LUT_B4F0 16'hB4C9
`define TANH_LUT_B4F8 16'hB4D1
`define TANH_LUT_B500 16'hB4D8
`define TANH_LUT_B508 16'hB4DF
`define TANH_LUT_B510 16'hB4E6
`define TANH_LUT_B518 16'hB4EE
`define TANH_LUT_B520 16'hB4F5
`define TANH_LUT_B528 16'hB4FC
`define TANH_LUT_B530 16'hB503
`define TANH_LUT_B538 16'hB50B
`define TANH_LUT_B540 16'hB512
`define TANH_LUT_B548 16'hB519
`define TANH_LUT_B550 16'hB520
`define TANH_LUT_B558 16'hB527
`define TANH_LUT_B560 16'hB52E
`define TANH_LUT_B568 16'hB536
`define TANH_LUT_B570 16'hB53D
`define TANH_LUT_B578 16'hB544
`define TANH_LUT_B580 16'hB54B
`define TANH_LUT_B588 16'hB552
`define TANH_LUT_B590 16'hB559
`define TANH_LUT_B598 16'hB560
`define TANH_LUT_B5A0 16'hB567
`define TANH_LUT_B5A8 16'hB56F
`define TANH_LUT_B5B0 16'hB576
`define TANH_LUT_B5B8 16'hB57D
`define TANH_LUT_B5C0 16'hB584
`define TANH_LUT_B5C8 16'hB58B
`define TANH_LUT_B5D0 16'hB592
`define TANH_LUT_B5D8 16'hB599
`define TANH_LUT_B5E0 16'hB5A0
`define TANH_LUT_B5E8 16'hB5A7
`define TANH_LUT_B5F0 16'hB5AE
`define TANH_LUT_B5F8 16'hB5B5
`define TANH_LUT_B600 16'hB5BC
`define TANH_LUT_B608 16'hB5C3
`define TANH_LUT_B610 16'hB5CA
`define TANH_LUT_B618 16'hB5D1
`define TANH_LUT_B620 16'hB5D8
`define TANH_LUT_B628 16'hB5DF
`define TANH_LUT_B630 16'hB5E5
`define TANH_LUT_B638 16'hB5EC
`define TANH_LUT_B640 16'hB5F3
`define TANH_LUT_B648 16'hB5FA
`define TANH_LUT_B650 16'hB601
`define TANH_LUT_B658 16'hB608
`define TANH_LUT_B660 16'hB60F
`define TANH_LUT_B668 16'hB616
`define TANH_LUT_B670 16'hB61C
`define TANH_LUT_B678 16'hB623
`define TANH_LUT_B680 16'hB62A
`define TANH_LUT_B688 16'hB631
`define TANH_LUT_B690 16'hB638
`define TANH_LUT_B698 16'hB63F
`define TANH_LUT_B6A0 16'hB645
`define TANH_LUT_B6A8 16'hB64C
`define TANH_LUT_B6B0 16'hB653
`define TANH_LUT_B6B8 16'hB65A
`define TANH_LUT_B6C0 16'hB660
`define TANH_LUT_B6C8 16'hB667
`define TANH_LUT_B6D0 16'hB66E
`define TANH_LUT_B6D8 16'hB674
`define TANH_LUT_B6E0 16'hB67B
`define TANH_LUT_B6E8 16'hB682
`define TANH_LUT_B6F0 16'hB688
`define TANH_LUT_B6F8 16'hB68F
`define TANH_LUT_B700 16'hB696
`define TANH_LUT_B708 16'hB69C
`define TANH_LUT_B710 16'hB6A3
`define TANH_LUT_B718 16'hB6AA
`define TANH_LUT_B720 16'hB6B0
`define TANH_LUT_B728 16'hB6B7
`define TANH_LUT_B730 16'hB6BD
`define TANH_LUT_B738 16'hB6C4
`define TANH_LUT_B740 16'hB6CB
`define TANH_LUT_B748 16'hB6D1
`define TANH_LUT_B750 16'hB6D8
`define TANH_LUT_B758 16'hB6DE
`define TANH_LUT_B760 16'hB6E5
`define TANH_LUT_B768 16'hB6EB
`define TANH_LUT_B770 16'hB6F2
`define TANH_LUT_B778 16'hB6F8
`define TANH_LUT_B780 16'hB6FF
`define TANH_LUT_B788 16'hB705
`define TANH_LUT_B790 16'hB70C
`define TANH_LUT_B798 16'hB712
`define TANH_LUT_B7A0 16'hB719
`define TANH_LUT_B7A8 16'hB71F
`define TANH_LUT_B7B0 16'hB725
`define TANH_LUT_B7B8 16'hB72C
`define TANH_LUT_B7C0 16'hB732
`define TANH_LUT_B7C8 16'hB739
`define TANH_LUT_B7D0 16'hB73F
`define TANH_LUT_B7D8 16'hB745
`define TANH_LUT_B7E0 16'hB74C
`define TANH_LUT_B7E8 16'hB752
`define TANH_LUT_B7F0 16'hB758
`define TANH_LUT_B7F8 16'hB75F
`define TANH_LUT_B800 16'hB765
`define TANH_LUT_B808 16'hB771
`define TANH_LUT_B810 16'hB77E
`define TANH_LUT_B818 16'hB78A
`define TANH_LUT_B820 16'hB797
`define TANH_LUT_B828 16'hB7A3
`define TANH_LUT_B830 16'hB7B0
`define TANH_LUT_B838 16'hB7BC
`define TANH_LUT_B840 16'hB7C8
`define TANH_LUT_B848 16'hB7D4
`define TANH_LUT_B850 16'hB7E0
`define TANH_LUT_B858 16'hB7EC
`define TANH_LUT_B860 16'hB7F9
`define TANH_LUT_B868 16'hB802
`define TANH_LUT_B870 16'hB808
`define TANH_LUT_B878 16'hB80E
`define TANH_LUT_B880 16'hB814
`define TANH_LUT_B888 16'hB81A
`define TANH_LUT_B890 16'hB820
`define TANH_LUT_B898 16'hB826
`define TANH_LUT_B8A0 16'hB82C
`define TANH_LUT_B8A8 16'hB831
`define TANH_LUT_B8B0 16'hB837
`define TANH_LUT_B8B8 16'hB83D
`define TANH_LUT_B8C0 16'hB843
`define TANH_LUT_B8C8 16'hB848
`define TANH_LUT_B8D0 16'hB84E
`define TANH_LUT_B8D8 16'hB854
`define TANH_LUT_B8E0 16'hB859
`define TANH_LUT_B8E8 16'hB85F
`define TANH_LUT_B8F0 16'hB865
`define TANH_LUT_B8F8 16'hB86A
`define TANH_LUT_B900 16'hB870
`define TANH_LUT_B908 16'hB875
`define TANH_LUT_B910 16'hB87B
`define TANH_LUT_B918 16'hB880
`define TANH_LUT_B920 16'hB886
`define TANH_LUT_B928 16'hB88B
`define TANH_LUT_B930 16'hB891
`define TANH_LUT_B938 16'hB896
`define TANH_LUT_B940 16'hB89B
`define TANH_LUT_B948 16'hB8A1
`define TANH_LUT_B950 16'hB8A6
`define TANH_LUT_B958 16'hB8AB
`define TANH_LUT_B960 16'hB8B1
`define TANH_LUT_B968 16'hB8B6
`define TANH_LUT_B970 16'hB8BB
`define TANH_LUT_B978 16'hB8C0
`define TANH_LUT_B980 16'hB8C5
`define TANH_LUT_B988 16'hB8CB
`define TANH_LUT_B990 16'hB8D0
`define TANH_LUT_B998 16'hB8D5
`define TANH_LUT_B9A0 16'hB8DA
`define TANH_LUT_B9A8 16'hB8DF
`define TANH_LUT_B9B0 16'hB8E4
`define TANH_LUT_B9B8 16'hB8E9
`define TANH_LUT_B9C0 16'hB8EE
`define TANH_LUT_B9C8 16'hB8F3
`define TANH_LUT_B9D0 16'hB8F8
`define TANH_LUT_B9D8 16'hB8FD
`define TANH_LUT_B9E0 16'hB902
`define TANH_LUT_B9E8 16'hB906
`define TANH_LUT_B9F0 16'hB90B
`define TANH_LUT_B9F8 16'hB910
`define TANH_LUT_BA00 16'hB915
`define TANH_LUT_BA08 16'hB91A
`define TANH_LUT_BA10 16'hB91E
`define TANH_LUT_BA18 16'hB923
`define TANH_LUT_BA20 16'hB928
`define TANH_LUT_BA28 16'hB92C
`define TANH_LUT_BA30 16'hB931
`define TANH_LUT_BA38 16'hB936
`define TANH_LUT_BA40 16'hB93A
`define TANH_LUT_BA48 16'hB93F
`define TANH_LUT_BA50 16'hB943
`define TANH_LUT_BA58 16'hB948
`define TANH_LUT_BA60 16'hB94C
`define TANH_LUT_BA68 16'hB951
`define TANH_LUT_BA70 16'hB955
`define TANH_LUT_BA78 16'hB95A
`define TANH_LUT_BA80 16'hB95E
`define TANH_LUT_BA88 16'hB963
`define TANH_LUT_BA90 16'hB967
`define TANH_LUT_BA98 16'hB96B
`define TANH_LUT_BAA0 16'hB970
`define TANH_LUT_BAA8 16'hB974
`define TANH_LUT_BAB0 16'hB978
`define TANH_LUT_BAB8 16'hB97C
`define TANH_LUT_BAC0 16'hB981
`define TANH_LUT_BAC8 16'hB985
`define TANH_LUT_BAD0 16'hB989
`define TANH_LUT_BAD8 16'hB98D
`define TANH_LUT_BAE0 16'hB991
`define TANH_LUT_BAE8 16'hB995
`define TANH_LUT_BAF0 16'hB999
`define TANH_LUT_BAF8 16'hB99E
`define TANH_LUT_BB00 16'hB9A2
`define TANH_LUT_BB08 16'hB9A6
`define TANH_LUT_BB10 16'hB9AA
`define TANH_LUT_BB18 16'hB9AE
`define TANH_LUT_BB20 16'hB9B2
`define TANH_LUT_BB28 16'hB9B6
`define TANH_LUT_BB30 16'hB9B9
`define TANH_LUT_BB38 16'hB9BD
`define TANH_LUT_BB40 16'hB9C1
`define TANH_LUT_BB48 16'hB9C5
`define TANH_LUT_BB50 16'hB9C9
`define TANH_LUT_BB58 16'hB9CD
`define TANH_LUT_BB60 16'hB9D0
`define TANH_LUT_BB68 16'hB9D4
`define TANH_LUT_BB70 16'hB9D8
`define TANH_LUT_BB78 16'hB9DC
`define TANH_LUT_BB80 16'hB9DF
`define TANH_LUT_BB88 16'hB9E3
`define TANH_LUT_BB90 16'hB9E7
`define TANH_LUT_BB98 16'hB9EA
`define TANH_LUT_BBA0 16'hB9EE
`define TANH_LUT_BBA8 16'hB9F2
`define TANH_LUT_BBB0 16'hB9F5
`define TANH_LUT_BBB8 16'hB9F9
`define TANH_LUT_BBC0 16'hB9FC
`define TANH_LUT_BBC8 16'hBA00
`define TANH_LUT_BBD0 16'hBA03
`define TANH_LUT_BBD8 16'hBA07
`define TANH_LUT_BBE0 16'hBA0A
`define TANH_LUT_BBE8 16'hBA0E
`define TANH_LUT_BBF0 16'hBA11
`define TANH_LUT_BBF8 16'hBA14
`define TANH_LUT_BC00 16'hBA18
`define TANH_LUT_BC08 16'hBA1E
`define TANH_LUT_BC10 16'hBA25
`define TANH_LUT_BC18 16'hBA2C
`define TANH_LUT_BC20 16'hBA32
`define TANH_LUT_BC28 16'hBA38
`define TANH_LUT_BC30 16'hBA3F
`define TANH_LUT_BC38 16'hBA45
`define TANH_LUT_BC40 16'hBA4B
`define TANH_LUT_BC48 16'hBA51
`define TANH_LUT_BC50 16'hBA57
`define TANH_LUT_BC58 16'hBA5D
`define TANH_LUT_BC60 16'hBA63
`define TANH_LUT_BC68 16'hBA69
`define TANH_LUT_BC70 16'hBA6E
`define TANH_LUT_BC78 16'hBA74
`define TANH_LUT_BC80 16'hBA79
`define TANH_LUT_BC88 16'hBA7F
`define TANH_LUT_BC90 16'hBA84
`define TANH_LUT_BC98 16'hBA8A
`define TANH_LUT_BCA0 16'hBA8F
`define TANH_LUT_BCA8 16'hBA94
`define TANH_LUT_BCB0 16'hBA99
`define TANH_LUT_BCB8 16'hBA9E
`define TANH_LUT_BCC0 16'hBAA3
`define TANH_LUT_BCC8 16'hBAA8
`define TANH_LUT_BCD0 16'hBAAD
`define TANH_LUT_BCD8 16'hBAB2
`define TANH_LUT_BCE0 16'hBAB7
`define TANH_LUT_BCE8 16'hBABC
`define TANH_LUT_BCF0 16'hBAC0
`define TANH_LUT_BCF8 16'hBAC5
`define TANH_LUT_BD00 16'hBAC9
`define TANH_LUT_BD08 16'hBACE
`define TANH_LUT_BD10 16'hBAD2
`define TANH_LUT_BD18 16'hBAD6
`define TANH_LUT_BD20 16'hBADB
`define TANH_LUT_BD28 16'hBADF
`define TANH_LUT_BD30 16'hBAE3
`define TANH_LUT_BD38 16'hBAE7
`define TANH_LUT_BD40 16'hBAEB
`define TANH_LUT_BD48 16'hBAEF
`define TANH_LUT_BD50 16'hBAF3
`define TANH_LUT_BD58 16'hBAF7
`define TANH_LUT_BD60 16'hBAFB
`define TANH_LUT_BD68 16'hBAFF
`define TANH_LUT_BD70 16'hBB03
`define TANH_LUT_BD78 16'hBB06
`define TANH_LUT_BD80 16'hBB0A
`define TANH_LUT_BD88 16'hBB0D
`define TANH_LUT_BD90 16'hBB11
`define TANH_LUT_BD98 16'hBB15
`define TANH_LUT_BDA0 16'hBB18
`define TANH_LUT_BDA8 16'hBB1B
`define TANH_LUT_BDB0 16'hBB1F
`define TANH_LUT_BDB8 16'hBB22
`define TANH_LUT_BDC0 16'hBB25
`define TANH_LUT_BDC8 16'hBB28
`define TANH_LUT_BDD0 16'hBB2C
`define TANH_LUT_BDD8 16'hBB2F
`define TANH_LUT_BDE0 16'hBB32
`define TANH_LUT_BDE8 16'hBB35
`define TANH_LUT_BDF0 16'hBB38
`define TANH_LUT_BDF8 16'hBB3B
`define TANH_LUT_BE00 16'hBB3E
`define TANH_LUT_BE08 16'hBB41
`define TANH_LUT_BE10 16'hBB43
`define TANH_LUT_BE18 16'hBB46
`define TANH_LUT_BE20 16'hBB49
`define TANH_LUT_BE28 16'hBB4C
`define TANH_LUT_BE30 16'hBB4E
`define TANH_LUT_BE38 16'hBB51
`define TANH_LUT_BE40 16'hBB54
`define TANH_LUT_BE48 16'hBB56
`define TANH_LUT_BE50 16'hBB59
`define TANH_LUT_BE58 16'hBB5B
`define TANH_LUT_BE60 16'hBB5E
`define TANH_LUT_BE68 16'hBB60
`define TANH_LUT_BE70 16'hBB62
`define TANH_LUT_BE78 16'hBB65
`define TANH_LUT_BE80 16'hBB67
`define TANH_LUT_BE88 16'hBB69
`define TANH_LUT_BE90 16'hBB6C
`define TANH_LUT_BE98 16'hBB6E
`define TANH_LUT_BEA0 16'hBB70
`define TANH_LUT_BEA8 16'hBB72
`define TANH_LUT_BEB0 16'hBB74
`define TANH_LUT_BEB8 16'hBB76
`define TANH_LUT_BEC0 16'hBB78
`define TANH_LUT_BEC8 16'hBB7B
`define TANH_LUT_BED0 16'hBB7D
`define TANH_LUT_BED8 16'hBB7E
`define TANH_LUT_BEE0 16'hBB80
`define TANH_LUT_BEE8 16'hBB82
`define TANH_LUT_BEF0 16'hBB84
`define TANH_LUT_BEF8 16'hBB86
`define TANH_LUT_BF00 16'hBB88
`define TANH_LUT_BF08 16'hBB8A
`define TANH_LUT_BF10 16'hBB8C
`define TANH_LUT_BF18 16'hBB8D
`define TANH_LUT_BF20 16'hBB8F
`define TANH_LUT_BF28 16'hBB91
`define TANH_LUT_BF30 16'hBB92
`define TANH_LUT_BF38 16'hBB94
`define TANH_LUT_BF40 16'hBB96
`define TANH_LUT_BF48 16'hBB97
`define TANH_LUT_BF50 16'hBB99
`define TANH_LUT_BF58 16'hBB9A
`define TANH_LUT_BF60 16'hBB9C
`define TANH_LUT_BF68 16'hBB9D
`define TANH_LUT_BF70 16'hBB9F
`define TANH_LUT_BF78 16'hBBA0
`define TANH_LUT_BF80 16'hBBA2
`define TANH_LUT_BF88 16'hBBA3
`define TANH_LUT_BF90 16'hBBA5
`define TANH_LUT_BF98 16'hBBA6
`define TANH_LUT_BFA0 16'hBBA7
`define TANH_LUT_BFA8 16'hBBA9
`define TANH_LUT_BFB0 16'hBBAA
`define TANH_LUT_BFB8 16'hBBAB
`define TANH_LUT_BFC0 16'hBBAD
`define TANH_LUT_BFC8 16'hBBAE
`define TANH_LUT_BFD0 16'hBBAF
`define TANH_LUT_BFD8 16'hBBB0
`define TANH_LUT_BFE0 16'hBBB2
`define TANH_LUT_BFE8 16'hBBB3
`define TANH_LUT_BFF0 16'hBBB4
`define TANH_LUT_BFF8 16'hBBB5
`define TANH_LUT_C000 16'hBBB6
`define TANH_LUT_C008 16'hBBB9
`define TANH_LUT_C010 16'hBBBB
`define TANH_LUT_C018 16'hBBBD
`define TANH_LUT_C020 16'hBBBF
`define TANH_LUT_C028 16'hBBC1
`define TANH_LUT_C030 16'hBBC3
`define TANH_LUT_C038 16'hBBC5
`define TANH_LUT_C040 16'hBBC6
`define TANH_LUT_C048 16'hBBC8
`define TANH_LUT_C050 16'hBBCA
`define TANH_LUT_C058 16'hBBCB
`define TANH_LUT_C060 16'hBBCD
`define TANH_LUT_C068 16'hBBCF
`define TANH_LUT_C070 16'hBBD0
`define TANH_LUT_C078 16'hBBD2
`define TANH_LUT_C080 16'hBBD3
`define TANH_LUT_C088 16'hBBD4
`define TANH_LUT_C090 16'hBBD6
`define TANH_LUT_C098 16'hBBD7
`define TANH_LUT_C0A0 16'hBBD8
`define TANH_LUT_C0A8 16'hBBD9
`define TANH_LUT_C0B0 16'hBBDB
`define TANH_LUT_C0B8 16'hBBDC
`define TANH_LUT_C0C0 16'hBBDD
`define TANH_LUT_C0C8 16'hBBDE
`define TANH_LUT_C0D0 16'hBBDF
`define TANH_LUT_C0D8 16'hBBE0
`define TANH_LUT_C0E0 16'hBBE1
`define TANH_LUT_C0E8 16'hBBE2
`define TANH_LUT_C0F0 16'hBBE3
`define TANH_LUT_C0F8 16'hBBE4
`define TANH_LUT_C100 16'hBBE5
`define TANH_LUT_C108 16'hBBE5
`define TANH_LUT_C110 16'hBBE6
`define TANH_LUT_C118 16'hBBE7
`define TANH_LUT_C120 16'hBBE8
`define TANH_LUT_C128 16'hBBE9
`define TANH_LUT_C130 16'hBBE9
`define TANH_LUT_C138 16'hBBEA
`define TANH_LUT_C140 16'hBBEB
`define TANH_LUT_C148 16'hBBEB
`define TANH_LUT_C150 16'hBBEC
`define TANH_LUT_C158 16'hBBED
`define TANH_LUT_C160 16'hBBED
`define TANH_LUT_C168 16'hBBEE
`define TANH_LUT_C170 16'hBBEE
`define TANH_LUT_C178 16'hBBEF
`define TANH_LUT_C180 16'hBBEF
`define TANH_LUT_C188 16'hBBF0
`define TANH_LUT_C190 16'hBBF0
`define TANH_LUT_C198 16'hBBF1
`define TANH_LUT_C1A0 16'hBBF1
`define TANH_LUT_C1A8 16'hBBF2
`define TANH_LUT_C1B0 16'hBBF2
`define TANH_LUT_C1B8 16'hBBF3
`define TANH_LUT_C1C0 16'hBBF3
`define TANH_LUT_C1C8 16'hBBF3
`define TANH_LUT_C1D0 16'hBBF4
`define TANH_LUT_C1D8 16'hBBF4
`define TANH_LUT_C1E0 16'hBBF5
`define TANH_LUT_C1E8 16'hBBF5
`define TANH_LUT_C1F0 16'hBBF5
`define TANH_LUT_C1F8 16'hBBF6
`define TANH_LUT_C200 16'hBBF6
`define TANH_LUT_C208 16'hBBF6
`define TANH_LUT_C210 16'hBBF6
`define TANH_LUT_C218 16'hBBF7
`define TANH_LUT_C220 16'hBBF7
`define TANH_LUT_C228 16'hBBF7
`define TANH_LUT_C230 16'hBBF8
`define TANH_LUT_C238 16'hBBF8
`define TANH_LUT_C240 16'hBBF8
`define TANH_LUT_C248 16'hBBF8
`define TANH_LUT_C250 16'hBBF9
`define TANH_LUT_C258 16'hBBF9
`define TANH_LUT_C260 16'hBBF9
`define TANH_LUT_C268 16'hBBF9
`define TANH_LUT_C270 16'hBBF9
`define TANH_LUT_C278 16'hBBFA
`define TANH_LUT_C280 16'hBBFA
`define TANH_LUT_C288 16'hBBFA
`define TANH_LUT_C290 16'hBBFA
`define TANH_LUT_C298 16'hBBFA
`define TANH_LUT_C2A0 16'hBBFB
`define TANH_LUT_C2A8 16'hBBFB
`define TANH_LUT_C2B0 16'hBBFB
`define TANH_LUT_C2B8 16'hBBFB
`define TANH_LUT_C2C0 16'hBBFB
`define TANH_LUT_C2C8 16'hBBFB
`define TANH_LUT_C2D0 16'hBBFB
`define TANH_LUT_C2D8 16'hBBFC
